module c6288 (N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528,N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288);
input N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528;
output N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288;
wire N546,N549,N552,N555,N558,N561,N564,N567,N570,N573,N576,N579,N582,N585,N588,N591,N594,N597,N600,N603,N606,N609,N612,N615,N618,N621,N624,N627,N630,N633,N636,N639,N642,N645,N648,N651,N654,N657,N660,N663,N666,N669,N672,N675,N678,N681,N684,N687,N690,N693,N696,N699,N702,N705,N708,N711,N714,N717,N720,N723,N726,N729,N732,N735,N738,N741,N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,N786,N789,N792,N795,N798,N801,N804,N807,N810,N813,N816,N819,N822,N825,N828,N831,N834,N837,N840,N843,N846,N849,N852,N855,N858,N861,N864,N867,N870,N873,N876,N879,N882,N885,N888,N891,N894,N897,N900,N903,N906,N909,N912,N915,N918,N921,N924,N927,N930,N933,N936,N939,N942,N945,N948,N951,N954,N957,N960,N963,N966,N969,N972,N975,N978,N981,N984,N987,N990,N993,N996,N999,N1002,N1005,N1008,N1011,N1014,N1017,N1020,N1023,N1026,N1029,N1032,N1035,N1038,N1041,N1044,N1047,N1050,N1053,N1056,N1059,N1062,N1065,N1068,N1071,N1074,N1077,N1080,N1083,N1086,N1089,N1092,N1095,N1098,N1101,N1104,N1107,N1110,N1113,N1116,N1119,N1122,N1125,N1128,N1131,N1134,N1137,N1140,N1143,N1146,N1149,N1152,N1155,N1158,N1161,N1164,N1167,N1170,N1173,N1176,N1179,N1182,N1185,N1188,N1191,N1194,N1197,N1200,N1203,N1206,N1209,N1212,N1215,N1218,N1221,N1224,N1227,N1230,N1233,N1236,N1239,N1242,N1245,N1248,N1251,N1254,N1257,N1260,N1263,N1266,N1269,N1272,N1275,N1278,N1281,N1284,N1287,N1290,N1293,N1296,N1299,N1302,N1305,N1308,N1311,N1315,N1319,N1323,N1327,N1331,N1335,N1339,N1343,N1347,N1351,N1355,N1359,N1363,N1367,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1450,N1454,N1458,N1462,N1466,N1470,N1474,N1478,N1482,N1486,N1490,N1494,N1498,N1502,N1506,N1507,N1508,N1511,N1512,N1513,N1516,N1517,N1518,N1521,N1522,N1523,N1526,N1527,N1528,N1531,N1532,N1533,N1536,N1537,N1538,N1541,N1542,N1543,N1546,N1547,N1548,N1551,N1552,N1553,N1556,N1557,N1558,N1561,N1562,N1563,N1566,N1567,N1568,N1571,N1572,N1573,N1576,N1577,N1578,N1582,N1585,N1588,N1591,N1594,N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,N1621,N1624,N1628,N1632,N1636,N1640,N1644,N1648,N1652,N1656,N1660,N1664,N1668,N1672,N1676,N1680,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1717,N1720,N1723,N1726,N1729,N1732,N1735,N1738,N1741,N1744,N1747,N1750,N1753,N1756,N1759,N1763,N1767,N1771,N1775,N1779,N1783,N1787,N1791,N1795,N1799,N1803,N1807,N1811,N1815,N1819,N1820,N1821,N1824,N1825,N1826,N1829,N1830,N1831,N1834,N1835,N1836,N1839,N1840,N1841,N1844,N1845,N1846,N1849,N1850,N1851,N1854,N1855,N1856,N1859,N1860,N1861,N1864,N1865,N1866,N1869,N1870,N1871,N1874,N1875,N1876,N1879,N1880,N1881,N1884,N1885,N1886,N1889,N1890,N1891,N1894,N1897,N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,N1932,N1935,N1938,N1941,N1945,N1946,N1947,N1951,N1955,N1959,N1963,N1967,N1971,N1975,N1979,N1983,N1987,N1991,N1995,N1999,N2000,N2001,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2033,N2037,N2040,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,N2067,N2070,N2073,N2076,N2080,N2081,N2082,N2085,N2089,N2093,N2097,N2101,N2105,N2109,N2113,N2117,N2121,N2125,N2129,N2133,N2137,N2138,N2139,N2142,N2145,N2149,N2150,N2151,N2154,N2155,N2156,N2159,N2160,N2161,N2164,N2165,N2166,N2169,N2170,N2171,N2174,N2175,N2176,N2179,N2180,N2181,N2184,N2185,N2186,N2189,N2190,N2191,N2194,N2195,N2196,N2199,N2200,N2201,N2204,N2205,N2206,N2209,N2210,N2211,N2214,N2217,N2221,N2222,N2224,N2227,N2230,N2233,N2236,N2239,N2242,N2245,N2248,N2251,N2254,N2257,N2260,N2264,N2265,N2266,N2269,N2273,N2277,N2281,N2285,N2289,N2293,N2297,N2301,N2305,N2309,N2313,N2317,N2318,N2319,N2322,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2353,N2357,N2358,N2359,N2362,N2365,N2368,N2371,N2374,N2377,N2380,N2383,N2386,N2389,N2392,N2395,N2398,N2402,N2403,N2404,N2407,N2410,N2414,N2418,N2422,N2426,N2430,N2434,N2438,N2442,N2446,N2450,N2454,N2458,N2462,N2463,N2464,N2467,N2470,N2474,N2475,N2476,N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2491,N2492,N2493,N2496,N2497,N2498,N2501,N2502,N2503,N2506,N2507,N2508,N2511,N2512,N2513,N2516,N2517,N2518,N2521,N2522,N2523,N2526,N2527,N2528,N2531,N2532,N2533,N2536,N2539,N2543,N2544,N2545,N2549,N2552,N2555,N2558,N2561,N2564,N2567,N2570,N2573,N2576,N2579,N2582,N2586,N2587,N2588,N2591,N2595,N2599,N2603,N2607,N2611,N2615,N2619,N2623,N2627,N2631,N2635,N2639,N2640,N2641,N2644,N2648,N2649,N2650,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2678,N2682,N2683,N2684,N2687,N2690,N2694,N2697,N2700,N2703,N2706,N2709,N2712,N2715,N2718,N2721,N2724,N2727,N2731,N2732,N2733,N2736,N2739,N2743,N2744,N2745,N2749,N2753,N2757,N2761,N2765,N2769,N2773,N2777,N2781,N2785,N2789,N2790,N2791,N2794,N2797,N2801,N2802,N2803,N2806,N2807,N2808,N2811,N2812,N2813,N2816,N2817,N2818,N2821,N2822,N2823,N2826,N2827,N2828,N2831,N2832,N2833,N2836,N2837,N2838,N2841,N2842,N2843,N2846,N2847,N2848,N2851,N2852,N2853,N2856,N2857,N2858,N2861,N2864,N2868,N2869,N2870,N2873,N2878,N2881,N2884,N2887,N2890,N2893,N2896,N2899,N2902,N2905,N2908,N2912,N2913,N2914,N2917,N2921,N2922,N2923,N2926,N2930,N2934,N2938,N2942,N2946,N2950,N2954,N2958,N2962,N2966,N2967,N2968,N2971,N2975,N2976,N2977,N2980,N2983,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3010,N3014,N3015,N3016,N3019,N3022,N3026,N3027,N3028,N3031,N3034,N3037,N3040,N3043,N3046,N3049,N3052,N3055,N3058,N3062,N3063,N3064,N3067,N3070,N3074,N3075,N3076,N3079,N3083,N3087,N3091,N3095,N3099,N3103,N3107,N3111,N3115,N3119,N3120,N3121,N3124,N3127,N3131,N3132,N3133,N3136,N3140,N3141,N3142,N3145,N3146,N3147,N3150,N3151,N3152,N3155,N3156,N3157,N3160,N3161,N3162,N3165,N3166,N3167,N3170,N3171,N3172,N3175,N3176,N3177,N3180,N3181,N3182,N3185,N3186,N3187,N3190,N3193,N3197,N3198,N3199,N3202,N3206,N3207,N3208,N3212,N3215,N3218,N3221,N3224,N3227,N3230,N3233,N3236,N3239,N3243,N3244,N3245,N3248,N3252,N3253,N3254,N3257,N3260,N3264,N3268,N3272,N3276,N3280,N3284,N3288,N3292,N3296,N3300,N3301,N3302,N3305,N3309,N3310,N3311,N3314,N3317,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3344,N3348,N3349,N3350,N3353,N3356,N3360,N3361,N3362,N3365,N3368,N3371,N3374,N3377,N3380,N3383,N3386,N3389,N3392,N3396,N3397,N3398,N3401,N3404,N3408,N3409,N3410,N3413,N3417,N3421,N3425,N3429,N3433,N3437,N3441,N3445,N3449,N3453,N3454,N3455,N3458,N3461,N3465,N3466,N3467,N3470,N3474,N3475,N3476,N3479,N3480,N3481,N3484,N3485,N3486,N3489,N3490,N3491,N3494,N3495,N3496,N3499,N3500,N3501,N3504,N3505,N3506,N3509,N3510,N3511,N3514,N3515,N3516,N3519,N3520,N3521,N3524,N3527,N3531,N3532,N3533,N3536,N3540,N3541,N3542,N3545,N3548,N3553,N3556,N3559,N3562,N3565,N3568,N3571,N3574,N3577,N3581,N3582,N3583,N3586,N3590,N3591,N3592,N3595,N3598,N3602,N3603,N3604,N3608,N3612,N3616,N3620,N3624,N3628,N3632,N3636,N3637,N3638,N3641,N3645,N3646,N3647,N3650,N3653,N3657,N3658,N3659,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3681,N3685,N3686,N3687,N3690,N3693,N3697,N3698,N3699,N3702,N3706,N3709,N3712,N3715,N3718,N3721,N3724,N3727,N3730,N3734,N3735,N3736,N3739,N3742,N3746,N3747,N3748,N3751,N3755,N3756,N3757,N3760,N3764,N3768,N3772,N3776,N3780,N3784,N3788,N3792,N3793,N3794,N3797,N3800,N3804,N3805,N3806,N3809,N3813,N3814,N3815,N3818,N3821,N3825,N3826,N3827,N3830,N3831,N3832,N3835,N3836,N3837,N3840,N3841,N3842,N3845,N3846,N3847,N3850,N3851,N3852,N3855,N3856,N3857,N3860,N3861,N3862,N3865,N3868,N3872,N3873,N3874,N3877,N3881,N3882,N3883,N3886,N3889,N3893,N3894,N3896,N3899,N3902,N3905,N3908,N3911,N3914,N3917,N3921,N3922,N3923,N3926,N3930,N3931,N3932,N3935,N3938,N3942,N3943,N3944,N3947,N3951,N3955,N3959,N3963,N3967,N3971,N3975,N3976,N3977,N3980,N3984,N3985,N3986,N3989,N3992,N3996,N3997,N3998,N4001,N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4022,N4026,N4027,N4028,N4031,N4034,N4038,N4039,N4040,N4043,N4047,N4048,N4049,N4052,N4055,N4058,N4061,N4064,N4067,N4070,N4073,N4077,N4078,N4079,N4082,N4085,N4089,N4090,N4091,N4094,N4098,N4099,N4100,N4103,N4106,N4110,N4114,N4118,N4122,N4126,N4130,N4134,N4138,N4139,N4140,N4143,N4146,N4150,N4151,N4152,N4155,N4159,N4160,N4161,N4164,N4167,N4171,N4172,N4173,N4174,N4175,N4178,N4179,N4180,N4183,N4184,N4185,N4188,N4189,N4190,N4193,N4194,N4195,N4198,N4199,N4200,N4203,N4204,N4205,N4208,N4211,N4215,N4216,N4217,N4220,N4224,N4225,N4226,N4229,N4232,N4236,N4237,N4238,N4242,N4245,N4248,N4251,N4254,N4257,N4260,N4264,N4265,N4266,N4269,N4273,N4274,N4275,N4278,N4281,N4285,N4286,N4287,N4290,N4294,N4298,N4302,N4306,N4310,N4314,N4318,N4319,N4320,N4323,N4327,N4328,N4329,N4332,N4335,N4339,N4340,N4341,N4344,N4348,N4349,N4350,N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4368,N4372,N4373,N4374,N4377,N4380,N4384,N4385,N4386,N4389,N4393,N4394,N4395,N4398,N4401,N4405,N4408,N4411,N4414,N4417,N4420,N4423,N4427,N4428,N4429,N4432,N4435,N4439,N4440,N4441,N4444,N4448,N4449,N4450,N4453,N4456,N4460,N4461,N4462,N4466,N4470,N4474,N4478,N4482,N4486,N4487,N4488,N4491,N4494,N4498,N4499,N4500,N4503,N4507,N4508,N4509,N4512,N4515,N4519,N4520,N4521,N4524,N4525,N4526,N4529,N4530,N4531,N4534,N4535,N4536,N4539,N4540,N4541,N4544,N4545,N4546,N4549,N4550,N4551,N4554,N4557,N4561,N4562,N4563,N4566,N4570,N4571,N4572,N4575,N4578,N4582,N4583,N4584,N4587,N4592,N4595,N4598,N4601,N4604,N4607,N4611,N4612,N4613,N4616,N4620,N4621,N4622,N4625,N4628,N4632,N4633,N4634,N4637,N4641,N4642,N4643,N4646,N4650,N4654,N4658,N4662,N4666,N4667,N4668,N4671,N4675,N4676,N4677,N4680,N4683,N4687,N4688,N4689,N4692,N4696,N4697,N4698,N4701,N4704,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718,N4721,N4725,N4726,N4727,N4730,N4733,N4737,N4738,N4739,N4742,N4746,N4747,N4748,N4751,N4754,N4758,N4759,N4760,N4763,N4766,N4769,N4772,N4775,N4779,N4780,N4781,N4784,N4787,N4791,N4792,N4793,N4796,N4800,N4801,N4802,N4805,N4808,N4812,N4813,N4814,N4817,N4821,N4825,N4829,N4833,N4837,N4838,N4839,N4842,N4845,N4849,N4850,N4851,N4854,N4858,N4859,N4860,N4863,N4866,N4870,N4871,N4872,N4875,N4879,N4880,N4881,N4884,N4885,N4886,N4889,N4890,N4891,N4894,N4895,N4896,N4899,N4900,N4901,N4904,N4907,N4911,N4912,N4913,N4916,N4920,N4921,N4922,N4925,N4928,N4932,N4933,N4934,N4937,N4941,N4942,N4943,N4947,N4950,N4953,N4956,N4959,N4963,N4964,N4965,N4968,N4972,N4973,N4974,N4977,N4980,N4984,N4985,N4986,N4989,N4993,N4994,N4995,N4998,N5001,N5005,N5009,N5013,N5017,N5021,N5022,N5023,N5026,N5030,N5031,N5032,N5035,N5038,N5042,N5043,N5044,N5047,N5051,N5052,N5053,N5056,N5059,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5076,N5080,N5081,N5082,N5085,N5088,N5092,N5093,N5094,N5097,N5101,N5102,N5103,N5106,N5109,N5113,N5114,N5115,N5118,N5121,N5124,N5127,N5130,N5134,N5135,N5136,N5139,N5142,N5146,N5147,N5148,N5151,N5155,N5156,N5157,N5160,N5163,N5167,N5168,N5169,N5172,N5176,N5180,N5184,N5188,N5192,N5193,N5194,N5197,N5200,N5204,N5205,N5206,N5209,N5213,N5214,N5215,N5218,N5221,N5225,N5226,N5227,N5230,N5234,N5235,N5236,N5239,N5240,N5241,N5244,N5245,N5246,N5249,N5250,N5251,N5254,N5255,N5256,N5259,N5262,N5266,N5267,N5268,N5271,N5275,N5276,N5277,N5280,N5283,N5287,N5288,N5289,N5292,N5296,N5297,N5298,N5301,N5304,N5309,N5312,N5315,N5318,N5322,N5323,N5324,N5327,N5331,N5332,N5333,N5336,N5339,N5343,N5344,N5345,N5348,N5352,N5353,N5354,N5357,N5360,N5364,N5365,N5366,N5370,N5374,N5378,N5379,N5380,N5383,N5387,N5388,N5389,N5392,N5395,N5399,N5400,N5401,N5404,N5408,N5409,N5410,N5413,N5416,N5420,N5421,N5422,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5434,N5438,N5439,N5440,N5443,N5446,N5450,N5451,N5452,N5455,N5459,N5460,N5461,N5464,N5467,N5471,N5472,N5473,N5476,N5480,N5483,N5486,N5489,N5493,N5494,N5495,N5498,N5501,N5505,N5506,N5507,N5510,N5514,N5515,N5516,N5519,N5522,N5526,N5527,N5528,N5531,N5535,N5536,N5537,N5540,N5544,N5548,N5552,N5553,N5554,N5557,N5560,N5564,N5565,N5566,N5569,N5573,N5574,N5575,N5578,N5581,N5585,N5586,N5587,N5590,N5594,N5595,N5596,N5599,N5602,N5606,N5607,N5608,N5611,N5612,N5613,N5616,N5617,N5618,N5621,N5624,N5628,N5629,N5630,N5633,N5637,N5638,N5639,N5642,N5645,N5649,N5650,N5651,N5654,N5658,N5659,N5660,N5663,N5666,N5670,N5671,N5673,N5676,N5679,N5683,N5684,N5685,N5688,N5692,N5693,N5694,N5697,N5700,N5704,N5705,N5706,N5709,N5713,N5714,N5715,N5718,N5721,N5725,N5726,N5727,N5730,N5734,N5738,N5739,N5740,N5743,N5747,N5748,N5749,N5752,N5755,N5759,N5760,N5761,N5764,N5768,N5769,N5770,N5773,N5776,N5780,N5781,N5782,N5785,N5786,N5787,N5788,N5789,N5792,N5796,N5797,N5798,N5801,N5804,N5808,N5809,N5810,N5813,N5817,N5818,N5819,N5822,N5825,N5829,N5830,N5831,N5834,N5837,N5840,N5844,N5845,N5846,N5849,N5852,N5856,N5857,N5858,N5861,N5865,N5866,N5867,N5870,N5873,N5877,N5878,N5879,N5882,N5886,N5890,N5891,N5892,N5895,N5898,N5902,N5903,N5904,N5907,N5911,N5912,N5913,N5916,N5919,N5923,N5924,N5925,N5928,N5929,N5930,N5933,N5934,N5935,N5938,N5941,N5945,N5946,N5947,N5950,N5954,N5955,N5956,N5959,N5962,N5966,N5967,N5968,N5972,N5975,N5979,N5980,N5981,N5984,N5988,N5989,N5990,N5993,N5996,N6000,N6001,N6002,N6005,N6009,N6010,N6011,N6014,N6018,N6019,N6020,N6023,N6026,N6030,N6031,N6032,N6035,N6036,N6037,N6040,N6044,N6045,N6046,N6049,N6052,N6056,N6057,N6058,N6061,N6064,N6068,N6069,N6070,N6073,N6076,N6080,N6081,N6082,N6085,N6089,N6090,N6091,N6094,N6097,N6101,N6102,N6103,N6106,N6107,N6108,N6111,N6114,N6118,N6119,N6120,N6124,N6128,N6129,N6130,N6133,N6134,N6135,N6138,N6141,N6145,N6146,N6147,N6151,N6155,N6156,N6157,N6161,N6165,N6166,N6167,N6171,N6175,N6176,N6177,N6181,N6185,N6186,N6187,N6191,N6195,N6196,N6197,N6201,N6205,N6206,N6207,N6211,N6215,N6216,N6217,N6221,N6225,N6226,N6227,N6231,N6235,N6236,N6237,N6241,N6245,N6246,N6247,N6251,N6255,N6256,N6257,N6261,N6265,N6266,N6267,N6271,N6275,N6276,N6277,N6281,N6285,N6286;
AND2X1 AND2_1 (.Y(N545),.A(N1),.B(N273));
AND2X1 AND2_2 (.Y(N546),.A(N1),.B(N290));
AND2X1 AND2_3 (.Y(N549),.A(N1),.B(N307));
AND2X1 AND2_4 (.Y(N552),.A(N1),.B(N324));
AND2X1 AND2_5 (.Y(N555),.A(N1),.B(N341));
AND2X1 AND2_6 (.Y(N558),.A(N1),.B(N358));
AND2X1 AND2_7 (.Y(N561),.A(N1),.B(N375));
AND2X1 AND2_8 (.Y(N564),.A(N1),.B(N392));
AND2X1 AND2_9 (.Y(N567),.A(N1),.B(N409));
AND2X1 AND2_10 (.Y(N570),.A(N1),.B(N426));
AND2X1 AND2_11 (.Y(N573),.A(N1),.B(N443));
AND2X1 AND2_12 (.Y(N576),.A(N1),.B(N460));
AND2X1 AND2_13 (.Y(N579),.A(N1),.B(N477));
AND2X1 AND2_14 (.Y(N582),.A(N1),.B(N494));
AND2X1 AND2_15 (.Y(N585),.A(N1),.B(N511));
AND2X1 AND2_16 (.Y(N588),.A(N1),.B(N528));
AND2X1 AND2_17 (.Y(N591),.A(N18),.B(N273));
AND2X1 AND2_18 (.Y(N594),.A(N18),.B(N290));
AND2X1 AND2_19 (.Y(N597),.A(N18),.B(N307));
AND2X1 AND2_20 (.Y(N600),.A(N18),.B(N324));
AND2X1 AND2_21 (.Y(N603),.A(N18),.B(N341));
AND2X1 AND2_22 (.Y(N606),.A(N18),.B(N358));
AND2X1 AND2_23 (.Y(N609),.A(N18),.B(N375));
AND2X1 AND2_24 (.Y(N612),.A(N18),.B(N392));
AND2X1 AND2_25 (.Y(N615),.A(N18),.B(N409));
AND2X1 AND2_26 (.Y(N618),.A(N18),.B(N426));
AND2X1 AND2_27 (.Y(N621),.A(N18),.B(N443));
AND2X1 AND2_28 (.Y(N624),.A(N18),.B(N460));
AND2X1 AND2_29 (.Y(N627),.A(N18),.B(N477));
AND2X1 AND2_30 (.Y(N630),.A(N18),.B(N494));
AND2X1 AND2_31 (.Y(N633),.A(N18),.B(N511));
AND2X1 AND2_32 (.Y(N636),.A(N18),.B(N528));
AND2X1 AND2_33 (.Y(N639),.A(N35),.B(N273));
AND2X1 AND2_34 (.Y(N642),.A(N35),.B(N290));
AND2X1 AND2_35 (.Y(N645),.A(N35),.B(N307));
AND2X1 AND2_36 (.Y(N648),.A(N35),.B(N324));
AND2X1 AND2_37 (.Y(N651),.A(N35),.B(N341));
AND2X1 AND2_38 (.Y(N654),.A(N35),.B(N358));
AND2X1 AND2_39 (.Y(N657),.A(N35),.B(N375));
AND2X1 AND2_40 (.Y(N660),.A(N35),.B(N392));
AND2X1 AND2_41 (.Y(N663),.A(N35),.B(N409));
AND2X1 AND2_42 (.Y(N666),.A(N35),.B(N426));
AND2X1 AND2_43 (.Y(N669),.A(N35),.B(N443));
AND2X1 AND2_44 (.Y(N672),.A(N35),.B(N460));
AND2X1 AND2_45 (.Y(N675),.A(N35),.B(N477));
AND2X1 AND2_46 (.Y(N678),.A(N35),.B(N494));
AND2X1 AND2_47 (.Y(N681),.A(N35),.B(N511));
AND2X1 AND2_48 (.Y(N684),.A(N35),.B(N528));
AND2X1 AND2_49 (.Y(N687),.A(N52),.B(N273));
AND2X1 AND2_50 (.Y(N690),.A(N52),.B(N290));
AND2X1 AND2_51 (.Y(N693),.A(N52),.B(N307));
AND2X1 AND2_52 (.Y(N696),.A(N52),.B(N324));
AND2X1 AND2_53 (.Y(N699),.A(N52),.B(N341));
AND2X1 AND2_54 (.Y(N702),.A(N52),.B(N358));
AND2X1 AND2_55 (.Y(N705),.A(N52),.B(N375));
AND2X1 AND2_56 (.Y(N708),.A(N52),.B(N392));
AND2X1 AND2_57 (.Y(N711),.A(N52),.B(N409));
AND2X1 AND2_58 (.Y(N714),.A(N52),.B(N426));
AND2X1 AND2_59 (.Y(N717),.A(N52),.B(N443));
AND2X1 AND2_60 (.Y(N720),.A(N52),.B(N460));
AND2X1 AND2_61 (.Y(N723),.A(N52),.B(N477));
AND2X1 AND2_62 (.Y(N726),.A(N52),.B(N494));
AND2X1 AND2_63 (.Y(N729),.A(N52),.B(N511));
AND2X1 AND2_64 (.Y(N732),.A(N52),.B(N528));
AND2X1 AND2_65 (.Y(N735),.A(N69),.B(N273));
AND2X1 AND2_66 (.Y(N738),.A(N69),.B(N290));
AND2X1 AND2_67 (.Y(N741),.A(N69),.B(N307));
AND2X1 AND2_68 (.Y(N744),.A(N69),.B(N324));
AND2X1 AND2_69 (.Y(N747),.A(N69),.B(N341));
AND2X1 AND2_70 (.Y(N750),.A(N69),.B(N358));
AND2X1 AND2_71 (.Y(N753),.A(N69),.B(N375));
AND2X1 AND2_72 (.Y(N756),.A(N69),.B(N392));
AND2X1 AND2_73 (.Y(N759),.A(N69),.B(N409));
AND2X1 AND2_74 (.Y(N762),.A(N69),.B(N426));
AND2X1 AND2_75 (.Y(N765),.A(N69),.B(N443));
AND2X1 AND2_76 (.Y(N768),.A(N69),.B(N460));
AND2X1 AND2_77 (.Y(N771),.A(N69),.B(N477));
AND2X1 AND2_78 (.Y(N774),.A(N69),.B(N494));
AND2X1 AND2_79 (.Y(N777),.A(N69),.B(N511));
AND2X1 AND2_80 (.Y(N780),.A(N69),.B(N528));
AND2X1 AND2_81 (.Y(N783),.A(N86),.B(N273));
AND2X1 AND2_82 (.Y(N786),.A(N86),.B(N290));
AND2X1 AND2_83 (.Y(N789),.A(N86),.B(N307));
AND2X1 AND2_84 (.Y(N792),.A(N86),.B(N324));
AND2X1 AND2_85 (.Y(N795),.A(N86),.B(N341));
AND2X1 AND2_86 (.Y(N798),.A(N86),.B(N358));
AND2X1 AND2_87 (.Y(N801),.A(N86),.B(N375));
AND2X1 AND2_88 (.Y(N804),.A(N86),.B(N392));
AND2X1 AND2_89 (.Y(N807),.A(N86),.B(N409));
AND2X1 AND2_90 (.Y(N810),.A(N86),.B(N426));
AND2X1 AND2_91 (.Y(N813),.A(N86),.B(N443));
AND2X1 AND2_92 (.Y(N816),.A(N86),.B(N460));
AND2X1 AND2_93 (.Y(N819),.A(N86),.B(N477));
AND2X1 AND2_94 (.Y(N822),.A(N86),.B(N494));
AND2X1 AND2_95 (.Y(N825),.A(N86),.B(N511));
AND2X1 AND2_96 (.Y(N828),.A(N86),.B(N528));
AND2X1 AND2_97 (.Y(N831),.A(N103),.B(N273));
AND2X1 AND2_98 (.Y(N834),.A(N103),.B(N290));
AND2X1 AND2_99 (.Y(N837),.A(N103),.B(N307));
AND2X1 AND2_100 (.Y(N840),.A(N103),.B(N324));
AND2X1 AND2_101 (.Y(N843),.A(N103),.B(N341));
AND2X1 AND2_102 (.Y(N846),.A(N103),.B(N358));
AND2X1 AND2_103 (.Y(N849),.A(N103),.B(N375));
AND2X1 AND2_104 (.Y(N852),.A(N103),.B(N392));
AND2X1 AND2_105 (.Y(N855),.A(N103),.B(N409));
AND2X1 AND2_106 (.Y(N858),.A(N103),.B(N426));
AND2X1 AND2_107 (.Y(N861),.A(N103),.B(N443));
AND2X1 AND2_108 (.Y(N864),.A(N103),.B(N460));
AND2X1 AND2_109 (.Y(N867),.A(N103),.B(N477));
AND2X1 AND2_110 (.Y(N870),.A(N103),.B(N494));
AND2X1 AND2_111 (.Y(N873),.A(N103),.B(N511));
AND2X1 AND2_112 (.Y(N876),.A(N103),.B(N528));
AND2X1 AND2_113 (.Y(N879),.A(N120),.B(N273));
AND2X1 AND2_114 (.Y(N882),.A(N120),.B(N290));
AND2X1 AND2_115 (.Y(N885),.A(N120),.B(N307));
AND2X1 AND2_116 (.Y(N888),.A(N120),.B(N324));
AND2X1 AND2_117 (.Y(N891),.A(N120),.B(N341));
AND2X1 AND2_118 (.Y(N894),.A(N120),.B(N358));
AND2X1 AND2_119 (.Y(N897),.A(N120),.B(N375));
AND2X1 AND2_120 (.Y(N900),.A(N120),.B(N392));
AND2X1 AND2_121 (.Y(N903),.A(N120),.B(N409));
AND2X1 AND2_122 (.Y(N906),.A(N120),.B(N426));
AND2X1 AND2_123 (.Y(N909),.A(N120),.B(N443));
AND2X1 AND2_124 (.Y(N912),.A(N120),.B(N460));
AND2X1 AND2_125 (.Y(N915),.A(N120),.B(N477));
AND2X1 AND2_126 (.Y(N918),.A(N120),.B(N494));
AND2X1 AND2_127 (.Y(N921),.A(N120),.B(N511));
AND2X1 AND2_128 (.Y(N924),.A(N120),.B(N528));
AND2X1 AND2_129 (.Y(N927),.A(N137),.B(N273));
AND2X1 AND2_130 (.Y(N930),.A(N137),.B(N290));
AND2X1 AND2_131 (.Y(N933),.A(N137),.B(N307));
AND2X1 AND2_132 (.Y(N936),.A(N137),.B(N324));
AND2X1 AND2_133 (.Y(N939),.A(N137),.B(N341));
AND2X1 AND2_134 (.Y(N942),.A(N137),.B(N358));
AND2X1 AND2_135 (.Y(N945),.A(N137),.B(N375));
AND2X1 AND2_136 (.Y(N948),.A(N137),.B(N392));
AND2X1 AND2_137 (.Y(N951),.A(N137),.B(N409));
AND2X1 AND2_138 (.Y(N954),.A(N137),.B(N426));
AND2X1 AND2_139 (.Y(N957),.A(N137),.B(N443));
AND2X1 AND2_140 (.Y(N960),.A(N137),.B(N460));
AND2X1 AND2_141 (.Y(N963),.A(N137),.B(N477));
AND2X1 AND2_142 (.Y(N966),.A(N137),.B(N494));
AND2X1 AND2_143 (.Y(N969),.A(N137),.B(N511));
AND2X1 AND2_144 (.Y(N972),.A(N137),.B(N528));
AND2X1 AND2_145 (.Y(N975),.A(N154),.B(N273));
AND2X1 AND2_146 (.Y(N978),.A(N154),.B(N290));
AND2X1 AND2_147 (.Y(N981),.A(N154),.B(N307));
AND2X1 AND2_148 (.Y(N984),.A(N154),.B(N324));
AND2X1 AND2_149 (.Y(N987),.A(N154),.B(N341));
AND2X1 AND2_150 (.Y(N990),.A(N154),.B(N358));
AND2X1 AND2_151 (.Y(N993),.A(N154),.B(N375));
AND2X1 AND2_152 (.Y(N996),.A(N154),.B(N392));
AND2X1 AND2_153 (.Y(N999),.A(N154),.B(N409));
AND2X1 AND2_154 (.Y(N1002),.A(N154),.B(N426));
AND2X1 AND2_155 (.Y(N1005),.A(N154),.B(N443));
AND2X1 AND2_156 (.Y(N1008),.A(N154),.B(N460));
AND2X1 AND2_157 (.Y(N1011),.A(N154),.B(N477));
AND2X1 AND2_158 (.Y(N1014),.A(N154),.B(N494));
AND2X1 AND2_159 (.Y(N1017),.A(N154),.B(N511));
AND2X1 AND2_160 (.Y(N1020),.A(N154),.B(N528));
AND2X1 AND2_161 (.Y(N1023),.A(N171),.B(N273));
AND2X1 AND2_162 (.Y(N1026),.A(N171),.B(N290));
AND2X1 AND2_163 (.Y(N1029),.A(N171),.B(N307));
AND2X1 AND2_164 (.Y(N1032),.A(N171),.B(N324));
AND2X1 AND2_165 (.Y(N1035),.A(N171),.B(N341));
AND2X1 AND2_166 (.Y(N1038),.A(N171),.B(N358));
AND2X1 AND2_167 (.Y(N1041),.A(N171),.B(N375));
AND2X1 AND2_168 (.Y(N1044),.A(N171),.B(N392));
AND2X1 AND2_169 (.Y(N1047),.A(N171),.B(N409));
AND2X1 AND2_170 (.Y(N1050),.A(N171),.B(N426));
AND2X1 AND2_171 (.Y(N1053),.A(N171),.B(N443));
AND2X1 AND2_172 (.Y(N1056),.A(N171),.B(N460));
AND2X1 AND2_173 (.Y(N1059),.A(N171),.B(N477));
AND2X1 AND2_174 (.Y(N1062),.A(N171),.B(N494));
AND2X1 AND2_175 (.Y(N1065),.A(N171),.B(N511));
AND2X1 AND2_176 (.Y(N1068),.A(N171),.B(N528));
AND2X1 AND2_177 (.Y(N1071),.A(N188),.B(N273));
AND2X1 AND2_178 (.Y(N1074),.A(N188),.B(N290));
AND2X1 AND2_179 (.Y(N1077),.A(N188),.B(N307));
AND2X1 AND2_180 (.Y(N1080),.A(N188),.B(N324));
AND2X1 AND2_181 (.Y(N1083),.A(N188),.B(N341));
AND2X1 AND2_182 (.Y(N1086),.A(N188),.B(N358));
AND2X1 AND2_183 (.Y(N1089),.A(N188),.B(N375));
AND2X1 AND2_184 (.Y(N1092),.A(N188),.B(N392));
AND2X1 AND2_185 (.Y(N1095),.A(N188),.B(N409));
AND2X1 AND2_186 (.Y(N1098),.A(N188),.B(N426));
AND2X1 AND2_187 (.Y(N1101),.A(N188),.B(N443));
AND2X1 AND2_188 (.Y(N1104),.A(N188),.B(N460));
AND2X1 AND2_189 (.Y(N1107),.A(N188),.B(N477));
AND2X1 AND2_190 (.Y(N1110),.A(N188),.B(N494));
AND2X1 AND2_191 (.Y(N1113),.A(N188),.B(N511));
AND2X1 AND2_192 (.Y(N1116),.A(N188),.B(N528));
AND2X1 AND2_193 (.Y(N1119),.A(N205),.B(N273));
AND2X1 AND2_194 (.Y(N1122),.A(N205),.B(N290));
AND2X1 AND2_195 (.Y(N1125),.A(N205),.B(N307));
AND2X1 AND2_196 (.Y(N1128),.A(N205),.B(N324));
AND2X1 AND2_197 (.Y(N1131),.A(N205),.B(N341));
AND2X1 AND2_198 (.Y(N1134),.A(N205),.B(N358));
AND2X1 AND2_199 (.Y(N1137),.A(N205),.B(N375));
AND2X1 AND2_200 (.Y(N1140),.A(N205),.B(N392));
AND2X1 AND2_201 (.Y(N1143),.A(N205),.B(N409));
AND2X1 AND2_202 (.Y(N1146),.A(N205),.B(N426));
AND2X1 AND2_203 (.Y(N1149),.A(N205),.B(N443));
AND2X1 AND2_204 (.Y(N1152),.A(N205),.B(N460));
AND2X1 AND2_205 (.Y(N1155),.A(N205),.B(N477));
AND2X1 AND2_206 (.Y(N1158),.A(N205),.B(N494));
AND2X1 AND2_207 (.Y(N1161),.A(N205),.B(N511));
AND2X1 AND2_208 (.Y(N1164),.A(N205),.B(N528));
AND2X1 AND2_209 (.Y(N1167),.A(N222),.B(N273));
AND2X1 AND2_210 (.Y(N1170),.A(N222),.B(N290));
AND2X1 AND2_211 (.Y(N1173),.A(N222),.B(N307));
AND2X1 AND2_212 (.Y(N1176),.A(N222),.B(N324));
AND2X1 AND2_213 (.Y(N1179),.A(N222),.B(N341));
AND2X1 AND2_214 (.Y(N1182),.A(N222),.B(N358));
AND2X1 AND2_215 (.Y(N1185),.A(N222),.B(N375));
AND2X1 AND2_216 (.Y(N1188),.A(N222),.B(N392));
AND2X1 AND2_217 (.Y(N1191),.A(N222),.B(N409));
AND2X1 AND2_218 (.Y(N1194),.A(N222),.B(N426));
AND2X1 AND2_219 (.Y(N1197),.A(N222),.B(N443));
AND2X1 AND2_220 (.Y(N1200),.A(N222),.B(N460));
AND2X1 AND2_221 (.Y(N1203),.A(N222),.B(N477));
AND2X1 AND2_222 (.Y(N1206),.A(N222),.B(N494));
AND2X1 AND2_223 (.Y(N1209),.A(N222),.B(N511));
AND2X1 AND2_224 (.Y(N1212),.A(N222),.B(N528));
AND2X1 AND2_225 (.Y(N1215),.A(N239),.B(N273));
AND2X1 AND2_226 (.Y(N1218),.A(N239),.B(N290));
AND2X1 AND2_227 (.Y(N1221),.A(N239),.B(N307));
AND2X1 AND2_228 (.Y(N1224),.A(N239),.B(N324));
AND2X1 AND2_229 (.Y(N1227),.A(N239),.B(N341));
AND2X1 AND2_230 (.Y(N1230),.A(N239),.B(N358));
AND2X1 AND2_231 (.Y(N1233),.A(N239),.B(N375));
AND2X1 AND2_232 (.Y(N1236),.A(N239),.B(N392));
AND2X1 AND2_233 (.Y(N1239),.A(N239),.B(N409));
AND2X1 AND2_234 (.Y(N1242),.A(N239),.B(N426));
AND2X1 AND2_235 (.Y(N1245),.A(N239),.B(N443));
AND2X1 AND2_236 (.Y(N1248),.A(N239),.B(N460));
AND2X1 AND2_237 (.Y(N1251),.A(N239),.B(N477));
AND2X1 AND2_238 (.Y(N1254),.A(N239),.B(N494));
AND2X1 AND2_239 (.Y(N1257),.A(N239),.B(N511));
AND2X1 AND2_240 (.Y(N1260),.A(N239),.B(N528));
AND2X1 AND2_241 (.Y(N1263),.A(N256),.B(N273));
AND2X1 AND2_242 (.Y(N1266),.A(N256),.B(N290));
AND2X1 AND2_243 (.Y(N1269),.A(N256),.B(N307));
AND2X1 AND2_244 (.Y(N1272),.A(N256),.B(N324));
AND2X1 AND2_245 (.Y(N1275),.A(N256),.B(N341));
AND2X1 AND2_246 (.Y(N1278),.A(N256),.B(N358));
AND2X1 AND2_247 (.Y(N1281),.A(N256),.B(N375));
AND2X1 AND2_248 (.Y(N1284),.A(N256),.B(N392));
AND2X1 AND2_249 (.Y(N1287),.A(N256),.B(N409));
AND2X1 AND2_250 (.Y(N1290),.A(N256),.B(N426));
AND2X1 AND2_251 (.Y(N1293),.A(N256),.B(N443));
AND2X1 AND2_252 (.Y(N1296),.A(N256),.B(N460));
AND2X1 AND2_253 (.Y(N1299),.A(N256),.B(N477));
AND2X1 AND2_254 (.Y(N1302),.A(N256),.B(N494));
AND2X1 AND2_255 (.Y(N1305),.A(N256),.B(N511));
AND2X1 AND2_256 (.Y(N1308),.A(N256),.B(N528));
INVX1 NOT1_257 (.Y(N1311),.A(N591));
INVX1 NOT1_258 (.Y(N1315),.A(N639));
INVX1 NOT1_259 (.Y(N1319),.A(N687));
INVX1 NOT1_260 (.Y(N1323),.A(N735));
INVX1 NOT1_261 (.Y(N1327),.A(N783));
INVX1 NOT1_262 (.Y(N1331),.A(N831));
INVX1 NOT1_263 (.Y(N1335),.A(N879));
INVX1 NOT1_264 (.Y(N1339),.A(N927));
INVX1 NOT1_265 (.Y(N1343),.A(N975));
INVX1 NOT1_266 (.Y(N1347),.A(N1023));
INVX1 NOT1_267 (.Y(N1351),.A(N1071));
INVX1 NOT1_268 (.Y(N1355),.A(N1119));
INVX1 NOT1_269 (.Y(N1359),.A(N1167));
INVX1 NOT1_270 (.Y(N1363),.A(N1215));
INVX1 NOT1_271 (.Y(N1367),.A(N1263));
NOR2X1 NOR2_272 (.Y(N1371),.A(N591),.B(N1311));
INVX1 NOT1_273 (.Y(N1372),.A(N1311));
NOR2X1 NOR2_274 (.Y(N1373),.A(N639),.B(N1315));
INVX1 NOT1_275 (.Y(N1374),.A(N1315));
NOR2X1 NOR2_276 (.Y(N1375),.A(N687),.B(N1319));
INVX1 NOT1_277 (.Y(N1376),.A(N1319));
NOR2X1 NOR2_278 (.Y(N1377),.A(N735),.B(N1323));
INVX1 NOT1_279 (.Y(N1378),.A(N1323));
NOR2X1 NOR2_280 (.Y(N1379),.A(N783),.B(N1327));
INVX1 NOT1_281 (.Y(N1380),.A(N1327));
NOR2X1 NOR2_282 (.Y(N1381),.A(N831),.B(N1331));
INVX1 NOT1_283 (.Y(N1382),.A(N1331));
NOR2X1 NOR2_284 (.Y(N1383),.A(N879),.B(N1335));
INVX1 NOT1_285 (.Y(N1384),.A(N1335));
NOR2X1 NOR2_286 (.Y(N1385),.A(N927),.B(N1339));
INVX1 NOT1_287 (.Y(N1386),.A(N1339));
NOR2X1 NOR2_288 (.Y(N1387),.A(N975),.B(N1343));
INVX1 NOT1_289 (.Y(N1388),.A(N1343));
NOR2X1 NOR2_290 (.Y(N1389),.A(N1023),.B(N1347));
INVX1 NOT1_291 (.Y(N1390),.A(N1347));
NOR2X1 NOR2_292 (.Y(N1391),.A(N1071),.B(N1351));
INVX1 NOT1_293 (.Y(N1392),.A(N1351));
NOR2X1 NOR2_294 (.Y(N1393),.A(N1119),.B(N1355));
INVX1 NOT1_295 (.Y(N1394),.A(N1355));
NOR2X1 NOR2_296 (.Y(N1395),.A(N1167),.B(N1359));
INVX1 NOT1_297 (.Y(N1396),.A(N1359));
NOR2X1 NOR2_298 (.Y(N1397),.A(N1215),.B(N1363));
INVX1 NOT1_299 (.Y(N1398),.A(N1363));
NOR2X1 NOR2_300 (.Y(N1399),.A(N1263),.B(N1367));
INVX1 NOT1_301 (.Y(N1400),.A(N1367));
NOR2X1 NOR2_302 (.Y(N1401),.A(N1371),.B(N1372));
NOR2X1 NOR2_303 (.Y(N1404),.A(N1373),.B(N1374));
NOR2X1 NOR2_304 (.Y(N1407),.A(N1375),.B(N1376));
NOR2X1 NOR2_305 (.Y(N1410),.A(N1377),.B(N1378));
NOR2X1 NOR2_306 (.Y(N1413),.A(N1379),.B(N1380));
NOR2X1 NOR2_307 (.Y(N1416),.A(N1381),.B(N1382));
NOR2X1 NOR2_308 (.Y(N1419),.A(N1383),.B(N1384));
NOR2X1 NOR2_309 (.Y(N1422),.A(N1385),.B(N1386));
NOR2X1 NOR2_310 (.Y(N1425),.A(N1387),.B(N1388));
NOR2X1 NOR2_311 (.Y(N1428),.A(N1389),.B(N1390));
NOR2X1 NOR2_312 (.Y(N1431),.A(N1391),.B(N1392));
NOR2X1 NOR2_313 (.Y(N1434),.A(N1393),.B(N1394));
NOR2X1 NOR2_314 (.Y(N1437),.A(N1395),.B(N1396));
NOR2X1 NOR2_315 (.Y(N1440),.A(N1397),.B(N1398));
NOR2X1 NOR2_316 (.Y(N1443),.A(N1399),.B(N1400));
NOR2X1 NOR2_317 (.Y(N1446),.A(N1401),.B(N546));
NOR2X1 NOR2_318 (.Y(N1450),.A(N1404),.B(N594));
NOR2X1 NOR2_319 (.Y(N1454),.A(N1407),.B(N642));
NOR2X1 NOR2_320 (.Y(N1458),.A(N1410),.B(N690));
NOR2X1 NOR2_321 (.Y(N1462),.A(N1413),.B(N738));
NOR2X1 NOR2_322 (.Y(N1466),.A(N1416),.B(N786));
NOR2X1 NOR2_323 (.Y(N1470),.A(N1419),.B(N834));
NOR2X1 NOR2_324 (.Y(N1474),.A(N1422),.B(N882));
NOR2X1 NOR2_325 (.Y(N1478),.A(N1425),.B(N930));
NOR2X1 NOR2_326 (.Y(N1482),.A(N1428),.B(N978));
NOR2X1 NOR2_327 (.Y(N1486),.A(N1431),.B(N1026));
NOR2X1 NOR2_328 (.Y(N1490),.A(N1434),.B(N1074));
NOR2X1 NOR2_329 (.Y(N1494),.A(N1437),.B(N1122));
NOR2X1 NOR2_330 (.Y(N1498),.A(N1440),.B(N1170));
NOR2X1 NOR2_331 (.Y(N1502),.A(N1443),.B(N1218));
NOR2X1 NOR2_332 (.Y(N1506),.A(N1401),.B(N1446));
NOR2X1 NOR2_333 (.Y(N1507),.A(N1446),.B(N546));
NOR2X1 NOR2_334 (.Y(N1508),.A(N1311),.B(N1446));
NOR2X1 NOR2_335 (.Y(N1511),.A(N1404),.B(N1450));
NOR2X1 NOR2_336 (.Y(N1512),.A(N1450),.B(N594));
NOR2X1 NOR2_337 (.Y(N1513),.A(N1315),.B(N1450));
NOR2X1 NOR2_338 (.Y(N1516),.A(N1407),.B(N1454));
NOR2X1 NOR2_339 (.Y(N1517),.A(N1454),.B(N642));
NOR2X1 NOR2_340 (.Y(N1518),.A(N1319),.B(N1454));
NOR2X1 NOR2_341 (.Y(N1521),.A(N1410),.B(N1458));
NOR2X1 NOR2_342 (.Y(N1522),.A(N1458),.B(N690));
NOR2X1 NOR2_343 (.Y(N1523),.A(N1323),.B(N1458));
NOR2X1 NOR2_344 (.Y(N1526),.A(N1413),.B(N1462));
NOR2X1 NOR2_345 (.Y(N1527),.A(N1462),.B(N738));
NOR2X1 NOR2_346 (.Y(N1528),.A(N1327),.B(N1462));
NOR2X1 NOR2_347 (.Y(N1531),.A(N1416),.B(N1466));
NOR2X1 NOR2_348 (.Y(N1532),.A(N1466),.B(N786));
NOR2X1 NOR2_349 (.Y(N1533),.A(N1331),.B(N1466));
NOR2X1 NOR2_350 (.Y(N1536),.A(N1419),.B(N1470));
NOR2X1 NOR2_351 (.Y(N1537),.A(N1470),.B(N834));
NOR2X1 NOR2_352 (.Y(N1538),.A(N1335),.B(N1470));
NOR2X1 NOR2_353 (.Y(N1541),.A(N1422),.B(N1474));
NOR2X1 NOR2_354 (.Y(N1542),.A(N1474),.B(N882));
NOR2X1 NOR2_355 (.Y(N1543),.A(N1339),.B(N1474));
NOR2X1 NOR2_356 (.Y(N1546),.A(N1425),.B(N1478));
NOR2X1 NOR2_357 (.Y(N1547),.A(N1478),.B(N930));
NOR2X1 NOR2_358 (.Y(N1548),.A(N1343),.B(N1478));
NOR2X1 NOR2_359 (.Y(N1551),.A(N1428),.B(N1482));
NOR2X1 NOR2_360 (.Y(N1552),.A(N1482),.B(N978));
NOR2X1 NOR2_361 (.Y(N1553),.A(N1347),.B(N1482));
NOR2X1 NOR2_362 (.Y(N1556),.A(N1431),.B(N1486));
NOR2X1 NOR2_363 (.Y(N1557),.A(N1486),.B(N1026));
NOR2X1 NOR2_364 (.Y(N1558),.A(N1351),.B(N1486));
NOR2X1 NOR2_365 (.Y(N1561),.A(N1434),.B(N1490));
NOR2X1 NOR2_366 (.Y(N1562),.A(N1490),.B(N1074));
NOR2X1 NOR2_367 (.Y(N1563),.A(N1355),.B(N1490));
NOR2X1 NOR2_368 (.Y(N1566),.A(N1437),.B(N1494));
NOR2X1 NOR2_369 (.Y(N1567),.A(N1494),.B(N1122));
NOR2X1 NOR2_370 (.Y(N1568),.A(N1359),.B(N1494));
NOR2X1 NOR2_371 (.Y(N1571),.A(N1440),.B(N1498));
NOR2X1 NOR2_372 (.Y(N1572),.A(N1498),.B(N1170));
NOR2X1 NOR2_373 (.Y(N1573),.A(N1363),.B(N1498));
NOR2X1 NOR2_374 (.Y(N1576),.A(N1443),.B(N1502));
NOR2X1 NOR2_375 (.Y(N1577),.A(N1502),.B(N1218));
NOR2X1 NOR2_376 (.Y(N1578),.A(N1367),.B(N1502));
NOR2X1 NOR2_377 (.Y(N1581),.A(N1506),.B(N1507));
NOR2X1 NOR2_378 (.Y(N1582),.A(N1511),.B(N1512));
NOR2X1 NOR2_379 (.Y(N1585),.A(N1516),.B(N1517));
NOR2X1 NOR2_380 (.Y(N1588),.A(N1521),.B(N1522));
NOR2X1 NOR2_381 (.Y(N1591),.A(N1526),.B(N1527));
NOR2X1 NOR2_382 (.Y(N1594),.A(N1531),.B(N1532));
NOR2X1 NOR2_383 (.Y(N1597),.A(N1536),.B(N1537));
NOR2X1 NOR2_384 (.Y(N1600),.A(N1541),.B(N1542));
NOR2X1 NOR2_385 (.Y(N1603),.A(N1546),.B(N1547));
NOR2X1 NOR2_386 (.Y(N1606),.A(N1551),.B(N1552));
NOR2X1 NOR2_387 (.Y(N1609),.A(N1556),.B(N1557));
NOR2X1 NOR2_388 (.Y(N1612),.A(N1561),.B(N1562));
NOR2X1 NOR2_389 (.Y(N1615),.A(N1566),.B(N1567));
NOR2X1 NOR2_390 (.Y(N1618),.A(N1571),.B(N1572));
NOR2X1 NOR2_391 (.Y(N1621),.A(N1576),.B(N1577));
NOR2X1 NOR2_392 (.Y(N1624),.A(N1266),.B(N1578));
NOR2X1 NOR2_393 (.Y(N1628),.A(N1582),.B(N1508));
NOR2X1 NOR2_394 (.Y(N1632),.A(N1585),.B(N1513));
NOR2X1 NOR2_395 (.Y(N1636),.A(N1588),.B(N1518));
NOR2X1 NOR2_396 (.Y(N1640),.A(N1591),.B(N1523));
NOR2X1 NOR2_397 (.Y(N1644),.A(N1594),.B(N1528));
NOR2X1 NOR2_398 (.Y(N1648),.A(N1597),.B(N1533));
NOR2X1 NOR2_399 (.Y(N1652),.A(N1600),.B(N1538));
NOR2X1 NOR2_400 (.Y(N1656),.A(N1603),.B(N1543));
NOR2X1 NOR2_401 (.Y(N1660),.A(N1606),.B(N1548));
NOR2X1 NOR2_402 (.Y(N1664),.A(N1609),.B(N1553));
NOR2X1 NOR2_403 (.Y(N1668),.A(N1612),.B(N1558));
NOR2X1 NOR2_404 (.Y(N1672),.A(N1615),.B(N1563));
NOR2X1 NOR2_405 (.Y(N1676),.A(N1618),.B(N1568));
NOR2X1 NOR2_406 (.Y(N1680),.A(N1621),.B(N1573));
NOR2X1 NOR2_407 (.Y(N1684),.A(N1266),.B(N1624));
NOR2X1 NOR2_408 (.Y(N1685),.A(N1624),.B(N1578));
NOR2X1 NOR2_409 (.Y(N1686),.A(N1582),.B(N1628));
NOR2X1 NOR2_410 (.Y(N1687),.A(N1628),.B(N1508));
NOR2X1 NOR2_411 (.Y(N1688),.A(N1585),.B(N1632));
NOR2X1 NOR2_412 (.Y(N1689),.A(N1632),.B(N1513));
NOR2X1 NOR2_413 (.Y(N1690),.A(N1588),.B(N1636));
NOR2X1 NOR2_414 (.Y(N1691),.A(N1636),.B(N1518));
NOR2X1 NOR2_415 (.Y(N1692),.A(N1591),.B(N1640));
NOR2X1 NOR2_416 (.Y(N1693),.A(N1640),.B(N1523));
NOR2X1 NOR2_417 (.Y(N1694),.A(N1594),.B(N1644));
NOR2X1 NOR2_418 (.Y(N1695),.A(N1644),.B(N1528));
NOR2X1 NOR2_419 (.Y(N1696),.A(N1597),.B(N1648));
NOR2X1 NOR2_420 (.Y(N1697),.A(N1648),.B(N1533));
NOR2X1 NOR2_421 (.Y(N1698),.A(N1600),.B(N1652));
NOR2X1 NOR2_422 (.Y(N1699),.A(N1652),.B(N1538));
NOR2X1 NOR2_423 (.Y(N1700),.A(N1603),.B(N1656));
NOR2X1 NOR2_424 (.Y(N1701),.A(N1656),.B(N1543));
NOR2X1 NOR2_425 (.Y(N1702),.A(N1606),.B(N1660));
NOR2X1 NOR2_426 (.Y(N1703),.A(N1660),.B(N1548));
NOR2X1 NOR2_427 (.Y(N1704),.A(N1609),.B(N1664));
NOR2X1 NOR2_428 (.Y(N1705),.A(N1664),.B(N1553));
NOR2X1 NOR2_429 (.Y(N1706),.A(N1612),.B(N1668));
NOR2X1 NOR2_430 (.Y(N1707),.A(N1668),.B(N1558));
NOR2X1 NOR2_431 (.Y(N1708),.A(N1615),.B(N1672));
NOR2X1 NOR2_432 (.Y(N1709),.A(N1672),.B(N1563));
NOR2X1 NOR2_433 (.Y(N1710),.A(N1618),.B(N1676));
NOR2X1 NOR2_434 (.Y(N1711),.A(N1676),.B(N1568));
NOR2X1 NOR2_435 (.Y(N1712),.A(N1621),.B(N1680));
NOR2X1 NOR2_436 (.Y(N1713),.A(N1680),.B(N1573));
NOR2X1 NOR2_437 (.Y(N1714),.A(N1684),.B(N1685));
NOR2X1 NOR2_438 (.Y(N1717),.A(N1686),.B(N1687));
NOR2X1 NOR2_439 (.Y(N1720),.A(N1688),.B(N1689));
NOR2X1 NOR2_440 (.Y(N1723),.A(N1690),.B(N1691));
NOR2X1 NOR2_441 (.Y(N1726),.A(N1692),.B(N1693));
NOR2X1 NOR2_442 (.Y(N1729),.A(N1694),.B(N1695));
NOR2X1 NOR2_443 (.Y(N1732),.A(N1696),.B(N1697));
NOR2X1 NOR2_444 (.Y(N1735),.A(N1698),.B(N1699));
NOR2X1 NOR2_445 (.Y(N1738),.A(N1700),.B(N1701));
NOR2X1 NOR2_446 (.Y(N1741),.A(N1702),.B(N1703));
NOR2X1 NOR2_447 (.Y(N1744),.A(N1704),.B(N1705));
NOR2X1 NOR2_448 (.Y(N1747),.A(N1706),.B(N1707));
NOR2X1 NOR2_449 (.Y(N1750),.A(N1708),.B(N1709));
NOR2X1 NOR2_450 (.Y(N1753),.A(N1710),.B(N1711));
NOR2X1 NOR2_451 (.Y(N1756),.A(N1712),.B(N1713));
NOR2X1 NOR2_452 (.Y(N1759),.A(N1714),.B(N1221));
NOR2X1 NOR2_453 (.Y(N1763),.A(N1717),.B(N549));
NOR2X1 NOR2_454 (.Y(N1767),.A(N1720),.B(N597));
NOR2X1 NOR2_455 (.Y(N1771),.A(N1723),.B(N645));
NOR2X1 NOR2_456 (.Y(N1775),.A(N1726),.B(N693));
NOR2X1 NOR2_457 (.Y(N1779),.A(N1729),.B(N741));
NOR2X1 NOR2_458 (.Y(N1783),.A(N1732),.B(N789));
NOR2X1 NOR2_459 (.Y(N1787),.A(N1735),.B(N837));
NOR2X1 NOR2_460 (.Y(N1791),.A(N1738),.B(N885));
NOR2X1 NOR2_461 (.Y(N1795),.A(N1741),.B(N933));
NOR2X1 NOR2_462 (.Y(N1799),.A(N1744),.B(N981));
NOR2X1 NOR2_463 (.Y(N1803),.A(N1747),.B(N1029));
NOR2X1 NOR2_464 (.Y(N1807),.A(N1750),.B(N1077));
NOR2X1 NOR2_465 (.Y(N1811),.A(N1753),.B(N1125));
NOR2X1 NOR2_466 (.Y(N1815),.A(N1756),.B(N1173));
NOR2X1 NOR2_467 (.Y(N1819),.A(N1714),.B(N1759));
NOR2X1 NOR2_468 (.Y(N1820),.A(N1759),.B(N1221));
NOR2X1 NOR2_469 (.Y(N1821),.A(N1624),.B(N1759));
NOR2X1 NOR2_470 (.Y(N1824),.A(N1717),.B(N1763));
NOR2X1 NOR2_471 (.Y(N1825),.A(N1763),.B(N549));
NOR2X1 NOR2_472 (.Y(N1826),.A(N1628),.B(N1763));
NOR2X1 NOR2_473 (.Y(N1829),.A(N1720),.B(N1767));
NOR2X1 NOR2_474 (.Y(N1830),.A(N1767),.B(N597));
NOR2X1 NOR2_475 (.Y(N1831),.A(N1632),.B(N1767));
NOR2X1 NOR2_476 (.Y(N1834),.A(N1723),.B(N1771));
NOR2X1 NOR2_477 (.Y(N1835),.A(N1771),.B(N645));
NOR2X1 NOR2_478 (.Y(N1836),.A(N1636),.B(N1771));
NOR2X1 NOR2_479 (.Y(N1839),.A(N1726),.B(N1775));
NOR2X1 NOR2_480 (.Y(N1840),.A(N1775),.B(N693));
NOR2X1 NOR2_481 (.Y(N1841),.A(N1640),.B(N1775));
NOR2X1 NOR2_482 (.Y(N1844),.A(N1729),.B(N1779));
NOR2X1 NOR2_483 (.Y(N1845),.A(N1779),.B(N741));
NOR2X1 NOR2_484 (.Y(N1846),.A(N1644),.B(N1779));
NOR2X1 NOR2_485 (.Y(N1849),.A(N1732),.B(N1783));
NOR2X1 NOR2_486 (.Y(N1850),.A(N1783),.B(N789));
NOR2X1 NOR2_487 (.Y(N1851),.A(N1648),.B(N1783));
NOR2X1 NOR2_488 (.Y(N1854),.A(N1735),.B(N1787));
NOR2X1 NOR2_489 (.Y(N1855),.A(N1787),.B(N837));
NOR2X1 NOR2_490 (.Y(N1856),.A(N1652),.B(N1787));
NOR2X1 NOR2_491 (.Y(N1859),.A(N1738),.B(N1791));
NOR2X1 NOR2_492 (.Y(N1860),.A(N1791),.B(N885));
NOR2X1 NOR2_493 (.Y(N1861),.A(N1656),.B(N1791));
NOR2X1 NOR2_494 (.Y(N1864),.A(N1741),.B(N1795));
NOR2X1 NOR2_495 (.Y(N1865),.A(N1795),.B(N933));
NOR2X1 NOR2_496 (.Y(N1866),.A(N1660),.B(N1795));
NOR2X1 NOR2_497 (.Y(N1869),.A(N1744),.B(N1799));
NOR2X1 NOR2_498 (.Y(N1870),.A(N1799),.B(N981));
NOR2X1 NOR2_499 (.Y(N1871),.A(N1664),.B(N1799));
NOR2X1 NOR2_500 (.Y(N1874),.A(N1747),.B(N1803));
NOR2X1 NOR2_501 (.Y(N1875),.A(N1803),.B(N1029));
NOR2X1 NOR2_502 (.Y(N1876),.A(N1668),.B(N1803));
NOR2X1 NOR2_503 (.Y(N1879),.A(N1750),.B(N1807));
NOR2X1 NOR2_504 (.Y(N1880),.A(N1807),.B(N1077));
NOR2X1 NOR2_505 (.Y(N1881),.A(N1672),.B(N1807));
NOR2X1 NOR2_506 (.Y(N1884),.A(N1753),.B(N1811));
NOR2X1 NOR2_507 (.Y(N1885),.A(N1811),.B(N1125));
NOR2X1 NOR2_508 (.Y(N1886),.A(N1676),.B(N1811));
NOR2X1 NOR2_509 (.Y(N1889),.A(N1756),.B(N1815));
NOR2X1 NOR2_510 (.Y(N1890),.A(N1815),.B(N1173));
NOR2X1 NOR2_511 (.Y(N1891),.A(N1680),.B(N1815));
NOR2X1 NOR2_512 (.Y(N1894),.A(N1819),.B(N1820));
NOR2X1 NOR2_513 (.Y(N1897),.A(N1269),.B(N1821));
NOR2X1 NOR2_514 (.Y(N1901),.A(N1824),.B(N1825));
NOR2X1 NOR2_515 (.Y(N1902),.A(N1829),.B(N1830));
NOR2X1 NOR2_516 (.Y(N1905),.A(N1834),.B(N1835));
NOR2X1 NOR2_517 (.Y(N1908),.A(N1839),.B(N1840));
NOR2X1 NOR2_518 (.Y(N1911),.A(N1844),.B(N1845));
NOR2X1 NOR2_519 (.Y(N1914),.A(N1849),.B(N1850));
NOR2X1 NOR2_520 (.Y(N1917),.A(N1854),.B(N1855));
NOR2X1 NOR2_521 (.Y(N1920),.A(N1859),.B(N1860));
NOR2X1 NOR2_522 (.Y(N1923),.A(N1864),.B(N1865));
NOR2X1 NOR2_523 (.Y(N1926),.A(N1869),.B(N1870));
NOR2X1 NOR2_524 (.Y(N1929),.A(N1874),.B(N1875));
NOR2X1 NOR2_525 (.Y(N1932),.A(N1879),.B(N1880));
NOR2X1 NOR2_526 (.Y(N1935),.A(N1884),.B(N1885));
NOR2X1 NOR2_527 (.Y(N1938),.A(N1889),.B(N1890));
NOR2X1 NOR2_528 (.Y(N1941),.A(N1894),.B(N1891));
NOR2X1 NOR2_529 (.Y(N1945),.A(N1269),.B(N1897));
NOR2X1 NOR2_530 (.Y(N1946),.A(N1897),.B(N1821));
NOR2X1 NOR2_531 (.Y(N1947),.A(N1902),.B(N1826));
NOR2X1 NOR2_532 (.Y(N1951),.A(N1905),.B(N1831));
NOR2X1 NOR2_533 (.Y(N1955),.A(N1908),.B(N1836));
NOR2X1 NOR2_534 (.Y(N1959),.A(N1911),.B(N1841));
NOR2X1 NOR2_535 (.Y(N1963),.A(N1914),.B(N1846));
NOR2X1 NOR2_536 (.Y(N1967),.A(N1917),.B(N1851));
NOR2X1 NOR2_537 (.Y(N1971),.A(N1920),.B(N1856));
NOR2X1 NOR2_538 (.Y(N1975),.A(N1923),.B(N1861));
NOR2X1 NOR2_539 (.Y(N1979),.A(N1926),.B(N1866));
NOR2X1 NOR2_540 (.Y(N1983),.A(N1929),.B(N1871));
NOR2X1 NOR2_541 (.Y(N1987),.A(N1932),.B(N1876));
NOR2X1 NOR2_542 (.Y(N1991),.A(N1935),.B(N1881));
NOR2X1 NOR2_543 (.Y(N1995),.A(N1938),.B(N1886));
NOR2X1 NOR2_544 (.Y(N1999),.A(N1894),.B(N1941));
NOR2X1 NOR2_545 (.Y(N2000),.A(N1941),.B(N1891));
NOR2X1 NOR2_546 (.Y(N2001),.A(N1945),.B(N1946));
NOR2X1 NOR2_547 (.Y(N2004),.A(N1902),.B(N1947));
NOR2X1 NOR2_548 (.Y(N2005),.A(N1947),.B(N1826));
NOR2X1 NOR2_549 (.Y(N2006),.A(N1905),.B(N1951));
NOR2X1 NOR2_550 (.Y(N2007),.A(N1951),.B(N1831));
NOR2X1 NOR2_551 (.Y(N2008),.A(N1908),.B(N1955));
NOR2X1 NOR2_552 (.Y(N2009),.A(N1955),.B(N1836));
NOR2X1 NOR2_553 (.Y(N2010),.A(N1911),.B(N1959));
NOR2X1 NOR2_554 (.Y(N2011),.A(N1959),.B(N1841));
NOR2X1 NOR2_555 (.Y(N2012),.A(N1914),.B(N1963));
NOR2X1 NOR2_556 (.Y(N2013),.A(N1963),.B(N1846));
NOR2X1 NOR2_557 (.Y(N2014),.A(N1917),.B(N1967));
NOR2X1 NOR2_558 (.Y(N2015),.A(N1967),.B(N1851));
NOR2X1 NOR2_559 (.Y(N2016),.A(N1920),.B(N1971));
NOR2X1 NOR2_560 (.Y(N2017),.A(N1971),.B(N1856));
NOR2X1 NOR2_561 (.Y(N2018),.A(N1923),.B(N1975));
NOR2X1 NOR2_562 (.Y(N2019),.A(N1975),.B(N1861));
NOR2X1 NOR2_563 (.Y(N2020),.A(N1926),.B(N1979));
NOR2X1 NOR2_564 (.Y(N2021),.A(N1979),.B(N1866));
NOR2X1 NOR2_565 (.Y(N2022),.A(N1929),.B(N1983));
NOR2X1 NOR2_566 (.Y(N2023),.A(N1983),.B(N1871));
NOR2X1 NOR2_567 (.Y(N2024),.A(N1932),.B(N1987));
NOR2X1 NOR2_568 (.Y(N2025),.A(N1987),.B(N1876));
NOR2X1 NOR2_569 (.Y(N2026),.A(N1935),.B(N1991));
NOR2X1 NOR2_570 (.Y(N2027),.A(N1991),.B(N1881));
NOR2X1 NOR2_571 (.Y(N2028),.A(N1938),.B(N1995));
NOR2X1 NOR2_572 (.Y(N2029),.A(N1995),.B(N1886));
NOR2X1 NOR2_573 (.Y(N2030),.A(N1999),.B(N2000));
NOR2X1 NOR2_574 (.Y(N2033),.A(N2001),.B(N1224));
NOR2X1 NOR2_575 (.Y(N2037),.A(N2004),.B(N2005));
NOR2X1 NOR2_576 (.Y(N2040),.A(N2006),.B(N2007));
NOR2X1 NOR2_577 (.Y(N2043),.A(N2008),.B(N2009));
NOR2X1 NOR2_578 (.Y(N2046),.A(N2010),.B(N2011));
NOR2X1 NOR2_579 (.Y(N2049),.A(N2012),.B(N2013));
NOR2X1 NOR2_580 (.Y(N2052),.A(N2014),.B(N2015));
NOR2X1 NOR2_581 (.Y(N2055),.A(N2016),.B(N2017));
NOR2X1 NOR2_582 (.Y(N2058),.A(N2018),.B(N2019));
NOR2X1 NOR2_583 (.Y(N2061),.A(N2020),.B(N2021));
NOR2X1 NOR2_584 (.Y(N2064),.A(N2022),.B(N2023));
NOR2X1 NOR2_585 (.Y(N2067),.A(N2024),.B(N2025));
NOR2X1 NOR2_586 (.Y(N2070),.A(N2026),.B(N2027));
NOR2X1 NOR2_587 (.Y(N2073),.A(N2028),.B(N2029));
NOR2X1 NOR2_588 (.Y(N2076),.A(N2030),.B(N1176));
NOR2X1 NOR2_589 (.Y(N2080),.A(N2001),.B(N2033));
NOR2X1 NOR2_590 (.Y(N2081),.A(N2033),.B(N1224));
NOR2X1 NOR2_591 (.Y(N2082),.A(N1897),.B(N2033));
NOR2X1 NOR2_592 (.Y(N2085),.A(N2037),.B(N552));
NOR2X1 NOR2_593 (.Y(N2089),.A(N2040),.B(N600));
NOR2X1 NOR2_594 (.Y(N2093),.A(N2043),.B(N648));
NOR2X1 NOR2_595 (.Y(N2097),.A(N2046),.B(N696));
NOR2X1 NOR2_596 (.Y(N2101),.A(N2049),.B(N744));
NOR2X1 NOR2_597 (.Y(N2105),.A(N2052),.B(N792));
NOR2X1 NOR2_598 (.Y(N2109),.A(N2055),.B(N840));
NOR2X1 NOR2_599 (.Y(N2113),.A(N2058),.B(N888));
NOR2X1 NOR2_600 (.Y(N2117),.A(N2061),.B(N936));
NOR2X1 NOR2_601 (.Y(N2121),.A(N2064),.B(N984));
NOR2X1 NOR2_602 (.Y(N2125),.A(N2067),.B(N1032));
NOR2X1 NOR2_603 (.Y(N2129),.A(N2070),.B(N1080));
NOR2X1 NOR2_604 (.Y(N2133),.A(N2073),.B(N1128));
NOR2X1 NOR2_605 (.Y(N2137),.A(N2030),.B(N2076));
NOR2X1 NOR2_606 (.Y(N2138),.A(N2076),.B(N1176));
NOR2X1 NOR2_607 (.Y(N2139),.A(N1941),.B(N2076));
NOR2X1 NOR2_608 (.Y(N2142),.A(N2080),.B(N2081));
NOR2X1 NOR2_609 (.Y(N2145),.A(N1272),.B(N2082));
NOR2X1 NOR2_610 (.Y(N2149),.A(N2037),.B(N2085));
NOR2X1 NOR2_611 (.Y(N2150),.A(N2085),.B(N552));
NOR2X1 NOR2_612 (.Y(N2151),.A(N1947),.B(N2085));
NOR2X1 NOR2_613 (.Y(N2154),.A(N2040),.B(N2089));
NOR2X1 NOR2_614 (.Y(N2155),.A(N2089),.B(N600));
NOR2X1 NOR2_615 (.Y(N2156),.A(N1951),.B(N2089));
NOR2X1 NOR2_616 (.Y(N2159),.A(N2043),.B(N2093));
NOR2X1 NOR2_617 (.Y(N2160),.A(N2093),.B(N648));
NOR2X1 NOR2_618 (.Y(N2161),.A(N1955),.B(N2093));
NOR2X1 NOR2_619 (.Y(N2164),.A(N2046),.B(N2097));
NOR2X1 NOR2_620 (.Y(N2165),.A(N2097),.B(N696));
NOR2X1 NOR2_621 (.Y(N2166),.A(N1959),.B(N2097));
NOR2X1 NOR2_622 (.Y(N2169),.A(N2049),.B(N2101));
NOR2X1 NOR2_623 (.Y(N2170),.A(N2101),.B(N744));
NOR2X1 NOR2_624 (.Y(N2171),.A(N1963),.B(N2101));
NOR2X1 NOR2_625 (.Y(N2174),.A(N2052),.B(N2105));
NOR2X1 NOR2_626 (.Y(N2175),.A(N2105),.B(N792));
NOR2X1 NOR2_627 (.Y(N2176),.A(N1967),.B(N2105));
NOR2X1 NOR2_628 (.Y(N2179),.A(N2055),.B(N2109));
NOR2X1 NOR2_629 (.Y(N2180),.A(N2109),.B(N840));
NOR2X1 NOR2_630 (.Y(N2181),.A(N1971),.B(N2109));
NOR2X1 NOR2_631 (.Y(N2184),.A(N2058),.B(N2113));
NOR2X1 NOR2_632 (.Y(N2185),.A(N2113),.B(N888));
NOR2X1 NOR2_633 (.Y(N2186),.A(N1975),.B(N2113));
NOR2X1 NOR2_634 (.Y(N2189),.A(N2061),.B(N2117));
NOR2X1 NOR2_635 (.Y(N2190),.A(N2117),.B(N936));
NOR2X1 NOR2_636 (.Y(N2191),.A(N1979),.B(N2117));
NOR2X1 NOR2_637 (.Y(N2194),.A(N2064),.B(N2121));
NOR2X1 NOR2_638 (.Y(N2195),.A(N2121),.B(N984));
NOR2X1 NOR2_639 (.Y(N2196),.A(N1983),.B(N2121));
NOR2X1 NOR2_640 (.Y(N2199),.A(N2067),.B(N2125));
NOR2X1 NOR2_641 (.Y(N2200),.A(N2125),.B(N1032));
NOR2X1 NOR2_642 (.Y(N2201),.A(N1987),.B(N2125));
NOR2X1 NOR2_643 (.Y(N2204),.A(N2070),.B(N2129));
NOR2X1 NOR2_644 (.Y(N2205),.A(N2129),.B(N1080));
NOR2X1 NOR2_645 (.Y(N2206),.A(N1991),.B(N2129));
NOR2X1 NOR2_646 (.Y(N2209),.A(N2073),.B(N2133));
NOR2X1 NOR2_647 (.Y(N2210),.A(N2133),.B(N1128));
NOR2X1 NOR2_648 (.Y(N2211),.A(N1995),.B(N2133));
NOR2X1 NOR2_649 (.Y(N2214),.A(N2137),.B(N2138));
NOR2X1 NOR2_650 (.Y(N2217),.A(N2142),.B(N2139));
NOR2X1 NOR2_651 (.Y(N2221),.A(N1272),.B(N2145));
NOR2X1 NOR2_652 (.Y(N2222),.A(N2145),.B(N2082));
NOR2X1 NOR2_653 (.Y(N2223),.A(N2149),.B(N2150));
NOR2X1 NOR2_654 (.Y(N2224),.A(N2154),.B(N2155));
NOR2X1 NOR2_655 (.Y(N2227),.A(N2159),.B(N2160));
NOR2X1 NOR2_656 (.Y(N2230),.A(N2164),.B(N2165));
NOR2X1 NOR2_657 (.Y(N2233),.A(N2169),.B(N2170));
NOR2X1 NOR2_658 (.Y(N2236),.A(N2174),.B(N2175));
NOR2X1 NOR2_659 (.Y(N2239),.A(N2179),.B(N2180));
NOR2X1 NOR2_660 (.Y(N2242),.A(N2184),.B(N2185));
NOR2X1 NOR2_661 (.Y(N2245),.A(N2189),.B(N2190));
NOR2X1 NOR2_662 (.Y(N2248),.A(N2194),.B(N2195));
NOR2X1 NOR2_663 (.Y(N2251),.A(N2199),.B(N2200));
NOR2X1 NOR2_664 (.Y(N2254),.A(N2204),.B(N2205));
NOR2X1 NOR2_665 (.Y(N2257),.A(N2209),.B(N2210));
NOR2X1 NOR2_666 (.Y(N2260),.A(N2214),.B(N2211));
NOR2X1 NOR2_667 (.Y(N2264),.A(N2142),.B(N2217));
NOR2X1 NOR2_668 (.Y(N2265),.A(N2217),.B(N2139));
NOR2X1 NOR2_669 (.Y(N2266),.A(N2221),.B(N2222));
NOR2X1 NOR2_670 (.Y(N2269),.A(N2224),.B(N2151));
NOR2X1 NOR2_671 (.Y(N2273),.A(N2227),.B(N2156));
NOR2X1 NOR2_672 (.Y(N2277),.A(N2230),.B(N2161));
NOR2X1 NOR2_673 (.Y(N2281),.A(N2233),.B(N2166));
NOR2X1 NOR2_674 (.Y(N2285),.A(N2236),.B(N2171));
NOR2X1 NOR2_675 (.Y(N2289),.A(N2239),.B(N2176));
NOR2X1 NOR2_676 (.Y(N2293),.A(N2242),.B(N2181));
NOR2X1 NOR2_677 (.Y(N2297),.A(N2245),.B(N2186));
NOR2X1 NOR2_678 (.Y(N2301),.A(N2248),.B(N2191));
NOR2X1 NOR2_679 (.Y(N2305),.A(N2251),.B(N2196));
NOR2X1 NOR2_680 (.Y(N2309),.A(N2254),.B(N2201));
NOR2X1 NOR2_681 (.Y(N2313),.A(N2257),.B(N2206));
NOR2X1 NOR2_682 (.Y(N2317),.A(N2214),.B(N2260));
NOR2X1 NOR2_683 (.Y(N2318),.A(N2260),.B(N2211));
NOR2X1 NOR2_684 (.Y(N2319),.A(N2264),.B(N2265));
NOR2X1 NOR2_685 (.Y(N2322),.A(N2266),.B(N1227));
NOR2X1 NOR2_686 (.Y(N2326),.A(N2224),.B(N2269));
NOR2X1 NOR2_687 (.Y(N2327),.A(N2269),.B(N2151));
NOR2X1 NOR2_688 (.Y(N2328),.A(N2227),.B(N2273));
NOR2X1 NOR2_689 (.Y(N2329),.A(N2273),.B(N2156));
NOR2X1 NOR2_690 (.Y(N2330),.A(N2230),.B(N2277));
NOR2X1 NOR2_691 (.Y(N2331),.A(N2277),.B(N2161));
NOR2X1 NOR2_692 (.Y(N2332),.A(N2233),.B(N2281));
NOR2X1 NOR2_693 (.Y(N2333),.A(N2281),.B(N2166));
NOR2X1 NOR2_694 (.Y(N2334),.A(N2236),.B(N2285));
NOR2X1 NOR2_695 (.Y(N2335),.A(N2285),.B(N2171));
NOR2X1 NOR2_696 (.Y(N2336),.A(N2239),.B(N2289));
NOR2X1 NOR2_697 (.Y(N2337),.A(N2289),.B(N2176));
NOR2X1 NOR2_698 (.Y(N2338),.A(N2242),.B(N2293));
NOR2X1 NOR2_699 (.Y(N2339),.A(N2293),.B(N2181));
NOR2X1 NOR2_700 (.Y(N2340),.A(N2245),.B(N2297));
NOR2X1 NOR2_701 (.Y(N2341),.A(N2297),.B(N2186));
NOR2X1 NOR2_702 (.Y(N2342),.A(N2248),.B(N2301));
NOR2X1 NOR2_703 (.Y(N2343),.A(N2301),.B(N2191));
NOR2X1 NOR2_704 (.Y(N2344),.A(N2251),.B(N2305));
NOR2X1 NOR2_705 (.Y(N2345),.A(N2305),.B(N2196));
NOR2X1 NOR2_706 (.Y(N2346),.A(N2254),.B(N2309));
NOR2X1 NOR2_707 (.Y(N2347),.A(N2309),.B(N2201));
NOR2X1 NOR2_708 (.Y(N2348),.A(N2257),.B(N2313));
NOR2X1 NOR2_709 (.Y(N2349),.A(N2313),.B(N2206));
NOR2X1 NOR2_710 (.Y(N2350),.A(N2317),.B(N2318));
NOR2X1 NOR2_711 (.Y(N2353),.A(N2319),.B(N1179));
NOR2X1 NOR2_712 (.Y(N2357),.A(N2266),.B(N2322));
NOR2X1 NOR2_713 (.Y(N2358),.A(N2322),.B(N1227));
NOR2X1 NOR2_714 (.Y(N2359),.A(N2145),.B(N2322));
NOR2X1 NOR2_715 (.Y(N2362),.A(N2326),.B(N2327));
NOR2X1 NOR2_716 (.Y(N2365),.A(N2328),.B(N2329));
NOR2X1 NOR2_717 (.Y(N2368),.A(N2330),.B(N2331));
NOR2X1 NOR2_718 (.Y(N2371),.A(N2332),.B(N2333));
NOR2X1 NOR2_719 (.Y(N2374),.A(N2334),.B(N2335));
NOR2X1 NOR2_720 (.Y(N2377),.A(N2336),.B(N2337));
NOR2X1 NOR2_721 (.Y(N2380),.A(N2338),.B(N2339));
NOR2X1 NOR2_722 (.Y(N2383),.A(N2340),.B(N2341));
NOR2X1 NOR2_723 (.Y(N2386),.A(N2342),.B(N2343));
NOR2X1 NOR2_724 (.Y(N2389),.A(N2344),.B(N2345));
NOR2X1 NOR2_725 (.Y(N2392),.A(N2346),.B(N2347));
NOR2X1 NOR2_726 (.Y(N2395),.A(N2348),.B(N2349));
NOR2X1 NOR2_727 (.Y(N2398),.A(N2350),.B(N1131));
NOR2X1 NOR2_728 (.Y(N2402),.A(N2319),.B(N2353));
NOR2X1 NOR2_729 (.Y(N2403),.A(N2353),.B(N1179));
NOR2X1 NOR2_730 (.Y(N2404),.A(N2217),.B(N2353));
NOR2X1 NOR2_731 (.Y(N2407),.A(N2357),.B(N2358));
NOR2X1 NOR2_732 (.Y(N2410),.A(N1275),.B(N2359));
NOR2X1 NOR2_733 (.Y(N2414),.A(N2362),.B(N555));
NOR2X1 NOR2_734 (.Y(N2418),.A(N2365),.B(N603));
NOR2X1 NOR2_735 (.Y(N2422),.A(N2368),.B(N651));
NOR2X1 NOR2_736 (.Y(N2426),.A(N2371),.B(N699));
NOR2X1 NOR2_737 (.Y(N2430),.A(N2374),.B(N747));
NOR2X1 NOR2_738 (.Y(N2434),.A(N2377),.B(N795));
NOR2X1 NOR2_739 (.Y(N2438),.A(N2380),.B(N843));
NOR2X1 NOR2_740 (.Y(N2442),.A(N2383),.B(N891));
NOR2X1 NOR2_741 (.Y(N2446),.A(N2386),.B(N939));
NOR2X1 NOR2_742 (.Y(N2450),.A(N2389),.B(N987));
NOR2X1 NOR2_743 (.Y(N2454),.A(N2392),.B(N1035));
NOR2X1 NOR2_744 (.Y(N2458),.A(N2395),.B(N1083));
NOR2X1 NOR2_745 (.Y(N2462),.A(N2350),.B(N2398));
NOR2X1 NOR2_746 (.Y(N2463),.A(N2398),.B(N1131));
NOR2X1 NOR2_747 (.Y(N2464),.A(N2260),.B(N2398));
NOR2X1 NOR2_748 (.Y(N2467),.A(N2402),.B(N2403));
NOR2X1 NOR2_749 (.Y(N2470),.A(N2407),.B(N2404));
NOR2X1 NOR2_750 (.Y(N2474),.A(N1275),.B(N2410));
NOR2X1 NOR2_751 (.Y(N2475),.A(N2410),.B(N2359));
NOR2X1 NOR2_752 (.Y(N2476),.A(N2362),.B(N2414));
NOR2X1 NOR2_753 (.Y(N2477),.A(N2414),.B(N555));
NOR2X1 NOR2_754 (.Y(N2478),.A(N2269),.B(N2414));
NOR2X1 NOR2_755 (.Y(N2481),.A(N2365),.B(N2418));
NOR2X1 NOR2_756 (.Y(N2482),.A(N2418),.B(N603));
NOR2X1 NOR2_757 (.Y(N2483),.A(N2273),.B(N2418));
NOR2X1 NOR2_758 (.Y(N2486),.A(N2368),.B(N2422));
NOR2X1 NOR2_759 (.Y(N2487),.A(N2422),.B(N651));
NOR2X1 NOR2_760 (.Y(N2488),.A(N2277),.B(N2422));
NOR2X1 NOR2_761 (.Y(N2491),.A(N2371),.B(N2426));
NOR2X1 NOR2_762 (.Y(N2492),.A(N2426),.B(N699));
NOR2X1 NOR2_763 (.Y(N2493),.A(N2281),.B(N2426));
NOR2X1 NOR2_764 (.Y(N2496),.A(N2374),.B(N2430));
NOR2X1 NOR2_765 (.Y(N2497),.A(N2430),.B(N747));
NOR2X1 NOR2_766 (.Y(N2498),.A(N2285),.B(N2430));
NOR2X1 NOR2_767 (.Y(N2501),.A(N2377),.B(N2434));
NOR2X1 NOR2_768 (.Y(N2502),.A(N2434),.B(N795));
NOR2X1 NOR2_769 (.Y(N2503),.A(N2289),.B(N2434));
NOR2X1 NOR2_770 (.Y(N2506),.A(N2380),.B(N2438));
NOR2X1 NOR2_771 (.Y(N2507),.A(N2438),.B(N843));
NOR2X1 NOR2_772 (.Y(N2508),.A(N2293),.B(N2438));
NOR2X1 NOR2_773 (.Y(N2511),.A(N2383),.B(N2442));
NOR2X1 NOR2_774 (.Y(N2512),.A(N2442),.B(N891));
NOR2X1 NOR2_775 (.Y(N2513),.A(N2297),.B(N2442));
NOR2X1 NOR2_776 (.Y(N2516),.A(N2386),.B(N2446));
NOR2X1 NOR2_777 (.Y(N2517),.A(N2446),.B(N939));
NOR2X1 NOR2_778 (.Y(N2518),.A(N2301),.B(N2446));
NOR2X1 NOR2_779 (.Y(N2521),.A(N2389),.B(N2450));
NOR2X1 NOR2_780 (.Y(N2522),.A(N2450),.B(N987));
NOR2X1 NOR2_781 (.Y(N2523),.A(N2305),.B(N2450));
NOR2X1 NOR2_782 (.Y(N2526),.A(N2392),.B(N2454));
NOR2X1 NOR2_783 (.Y(N2527),.A(N2454),.B(N1035));
NOR2X1 NOR2_784 (.Y(N2528),.A(N2309),.B(N2454));
NOR2X1 NOR2_785 (.Y(N2531),.A(N2395),.B(N2458));
NOR2X1 NOR2_786 (.Y(N2532),.A(N2458),.B(N1083));
NOR2X1 NOR2_787 (.Y(N2533),.A(N2313),.B(N2458));
NOR2X1 NOR2_788 (.Y(N2536),.A(N2462),.B(N2463));
NOR2X1 NOR2_789 (.Y(N2539),.A(N2467),.B(N2464));
NOR2X1 NOR2_790 (.Y(N2543),.A(N2407),.B(N2470));
NOR2X1 NOR2_791 (.Y(N2544),.A(N2470),.B(N2404));
NOR2X1 NOR2_792 (.Y(N2545),.A(N2474),.B(N2475));
NOR2X1 NOR2_793 (.Y(N2548),.A(N2476),.B(N2477));
NOR2X1 NOR2_794 (.Y(N2549),.A(N2481),.B(N2482));
NOR2X1 NOR2_795 (.Y(N2552),.A(N2486),.B(N2487));
NOR2X1 NOR2_796 (.Y(N2555),.A(N2491),.B(N2492));
NOR2X1 NOR2_797 (.Y(N2558),.A(N2496),.B(N2497));
NOR2X1 NOR2_798 (.Y(N2561),.A(N2501),.B(N2502));
NOR2X1 NOR2_799 (.Y(N2564),.A(N2506),.B(N2507));
NOR2X1 NOR2_800 (.Y(N2567),.A(N2511),.B(N2512));
NOR2X1 NOR2_801 (.Y(N2570),.A(N2516),.B(N2517));
NOR2X1 NOR2_802 (.Y(N2573),.A(N2521),.B(N2522));
NOR2X1 NOR2_803 (.Y(N2576),.A(N2526),.B(N2527));
NOR2X1 NOR2_804 (.Y(N2579),.A(N2531),.B(N2532));
NOR2X1 NOR2_805 (.Y(N2582),.A(N2536),.B(N2533));
NOR2X1 NOR2_806 (.Y(N2586),.A(N2467),.B(N2539));
NOR2X1 NOR2_807 (.Y(N2587),.A(N2539),.B(N2464));
NOR2X1 NOR2_808 (.Y(N2588),.A(N2543),.B(N2544));
NOR2X1 NOR2_809 (.Y(N2591),.A(N2545),.B(N1230));
NOR2X1 NOR2_810 (.Y(N2595),.A(N2549),.B(N2478));
NOR2X1 NOR2_811 (.Y(N2599),.A(N2552),.B(N2483));
NOR2X1 NOR2_812 (.Y(N2603),.A(N2555),.B(N2488));
NOR2X1 NOR2_813 (.Y(N2607),.A(N2558),.B(N2493));
NOR2X1 NOR2_814 (.Y(N2611),.A(N2561),.B(N2498));
NOR2X1 NOR2_815 (.Y(N2615),.A(N2564),.B(N2503));
NOR2X1 NOR2_816 (.Y(N2619),.A(N2567),.B(N2508));
NOR2X1 NOR2_817 (.Y(N2623),.A(N2570),.B(N2513));
NOR2X1 NOR2_818 (.Y(N2627),.A(N2573),.B(N2518));
NOR2X1 NOR2_819 (.Y(N2631),.A(N2576),.B(N2523));
NOR2X1 NOR2_820 (.Y(N2635),.A(N2579),.B(N2528));
NOR2X1 NOR2_821 (.Y(N2639),.A(N2536),.B(N2582));
NOR2X1 NOR2_822 (.Y(N2640),.A(N2582),.B(N2533));
NOR2X1 NOR2_823 (.Y(N2641),.A(N2586),.B(N2587));
NOR2X1 NOR2_824 (.Y(N2644),.A(N2588),.B(N1182));
NOR2X1 NOR2_825 (.Y(N2648),.A(N2545),.B(N2591));
NOR2X1 NOR2_826 (.Y(N2649),.A(N2591),.B(N1230));
NOR2X1 NOR2_827 (.Y(N2650),.A(N2410),.B(N2591));
NOR2X1 NOR2_828 (.Y(N2653),.A(N2549),.B(N2595));
NOR2X1 NOR2_829 (.Y(N2654),.A(N2595),.B(N2478));
NOR2X1 NOR2_830 (.Y(N2655),.A(N2552),.B(N2599));
NOR2X1 NOR2_831 (.Y(N2656),.A(N2599),.B(N2483));
NOR2X1 NOR2_832 (.Y(N2657),.A(N2555),.B(N2603));
NOR2X1 NOR2_833 (.Y(N2658),.A(N2603),.B(N2488));
NOR2X1 NOR2_834 (.Y(N2659),.A(N2558),.B(N2607));
NOR2X1 NOR2_835 (.Y(N2660),.A(N2607),.B(N2493));
NOR2X1 NOR2_836 (.Y(N2661),.A(N2561),.B(N2611));
NOR2X1 NOR2_837 (.Y(N2662),.A(N2611),.B(N2498));
NOR2X1 NOR2_838 (.Y(N2663),.A(N2564),.B(N2615));
NOR2X1 NOR2_839 (.Y(N2664),.A(N2615),.B(N2503));
NOR2X1 NOR2_840 (.Y(N2665),.A(N2567),.B(N2619));
NOR2X1 NOR2_841 (.Y(N2666),.A(N2619),.B(N2508));
NOR2X1 NOR2_842 (.Y(N2667),.A(N2570),.B(N2623));
NOR2X1 NOR2_843 (.Y(N2668),.A(N2623),.B(N2513));
NOR2X1 NOR2_844 (.Y(N2669),.A(N2573),.B(N2627));
NOR2X1 NOR2_845 (.Y(N2670),.A(N2627),.B(N2518));
NOR2X1 NOR2_846 (.Y(N2671),.A(N2576),.B(N2631));
NOR2X1 NOR2_847 (.Y(N2672),.A(N2631),.B(N2523));
NOR2X1 NOR2_848 (.Y(N2673),.A(N2579),.B(N2635));
NOR2X1 NOR2_849 (.Y(N2674),.A(N2635),.B(N2528));
NOR2X1 NOR2_850 (.Y(N2675),.A(N2639),.B(N2640));
NOR2X1 NOR2_851 (.Y(N2678),.A(N2641),.B(N1134));
NOR2X1 NOR2_852 (.Y(N2682),.A(N2588),.B(N2644));
NOR2X1 NOR2_853 (.Y(N2683),.A(N2644),.B(N1182));
NOR2X1 NOR2_854 (.Y(N2684),.A(N2470),.B(N2644));
NOR2X1 NOR2_855 (.Y(N2687),.A(N2648),.B(N2649));
NOR2X1 NOR2_856 (.Y(N2690),.A(N1278),.B(N2650));
NOR2X1 NOR2_857 (.Y(N2694),.A(N2653),.B(N2654));
NOR2X1 NOR2_858 (.Y(N2697),.A(N2655),.B(N2656));
NOR2X1 NOR2_859 (.Y(N2700),.A(N2657),.B(N2658));
NOR2X1 NOR2_860 (.Y(N2703),.A(N2659),.B(N2660));
NOR2X1 NOR2_861 (.Y(N2706),.A(N2661),.B(N2662));
NOR2X1 NOR2_862 (.Y(N2709),.A(N2663),.B(N2664));
NOR2X1 NOR2_863 (.Y(N2712),.A(N2665),.B(N2666));
NOR2X1 NOR2_864 (.Y(N2715),.A(N2667),.B(N2668));
NOR2X1 NOR2_865 (.Y(N2718),.A(N2669),.B(N2670));
NOR2X1 NOR2_866 (.Y(N2721),.A(N2671),.B(N2672));
NOR2X1 NOR2_867 (.Y(N2724),.A(N2673),.B(N2674));
NOR2X1 NOR2_868 (.Y(N2727),.A(N2675),.B(N1086));
NOR2X1 NOR2_869 (.Y(N2731),.A(N2641),.B(N2678));
NOR2X1 NOR2_870 (.Y(N2732),.A(N2678),.B(N1134));
NOR2X1 NOR2_871 (.Y(N2733),.A(N2539),.B(N2678));
NOR2X1 NOR2_872 (.Y(N2736),.A(N2682),.B(N2683));
NOR2X1 NOR2_873 (.Y(N2739),.A(N2687),.B(N2684));
NOR2X1 NOR2_874 (.Y(N2743),.A(N1278),.B(N2690));
NOR2X1 NOR2_875 (.Y(N2744),.A(N2690),.B(N2650));
NOR2X1 NOR2_876 (.Y(N2745),.A(N2694),.B(N558));
NOR2X1 NOR2_877 (.Y(N2749),.A(N2697),.B(N606));
NOR2X1 NOR2_878 (.Y(N2753),.A(N2700),.B(N654));
NOR2X1 NOR2_879 (.Y(N2757),.A(N2703),.B(N702));
NOR2X1 NOR2_880 (.Y(N2761),.A(N2706),.B(N750));
NOR2X1 NOR2_881 (.Y(N2765),.A(N2709),.B(N798));
NOR2X1 NOR2_882 (.Y(N2769),.A(N2712),.B(N846));
NOR2X1 NOR2_883 (.Y(N2773),.A(N2715),.B(N894));
NOR2X1 NOR2_884 (.Y(N2777),.A(N2718),.B(N942));
NOR2X1 NOR2_885 (.Y(N2781),.A(N2721),.B(N990));
NOR2X1 NOR2_886 (.Y(N2785),.A(N2724),.B(N1038));
NOR2X1 NOR2_887 (.Y(N2789),.A(N2675),.B(N2727));
NOR2X1 NOR2_888 (.Y(N2790),.A(N2727),.B(N1086));
NOR2X1 NOR2_889 (.Y(N2791),.A(N2582),.B(N2727));
NOR2X1 NOR2_890 (.Y(N2794),.A(N2731),.B(N2732));
NOR2X1 NOR2_891 (.Y(N2797),.A(N2736),.B(N2733));
NOR2X1 NOR2_892 (.Y(N2801),.A(N2687),.B(N2739));
NOR2X1 NOR2_893 (.Y(N2802),.A(N2739),.B(N2684));
NOR2X1 NOR2_894 (.Y(N2803),.A(N2743),.B(N2744));
NOR2X1 NOR2_895 (.Y(N2806),.A(N2694),.B(N2745));
NOR2X1 NOR2_896 (.Y(N2807),.A(N2745),.B(N558));
NOR2X1 NOR2_897 (.Y(N2808),.A(N2595),.B(N2745));
NOR2X1 NOR2_898 (.Y(N2811),.A(N2697),.B(N2749));
NOR2X1 NOR2_899 (.Y(N2812),.A(N2749),.B(N606));
NOR2X1 NOR2_900 (.Y(N2813),.A(N2599),.B(N2749));
NOR2X1 NOR2_901 (.Y(N2816),.A(N2700),.B(N2753));
NOR2X1 NOR2_902 (.Y(N2817),.A(N2753),.B(N654));
NOR2X1 NOR2_903 (.Y(N2818),.A(N2603),.B(N2753));
NOR2X1 NOR2_904 (.Y(N2821),.A(N2703),.B(N2757));
NOR2X1 NOR2_905 (.Y(N2822),.A(N2757),.B(N702));
NOR2X1 NOR2_906 (.Y(N2823),.A(N2607),.B(N2757));
NOR2X1 NOR2_907 (.Y(N2826),.A(N2706),.B(N2761));
NOR2X1 NOR2_908 (.Y(N2827),.A(N2761),.B(N750));
NOR2X1 NOR2_909 (.Y(N2828),.A(N2611),.B(N2761));
NOR2X1 NOR2_910 (.Y(N2831),.A(N2709),.B(N2765));
NOR2X1 NOR2_911 (.Y(N2832),.A(N2765),.B(N798));
NOR2X1 NOR2_912 (.Y(N2833),.A(N2615),.B(N2765));
NOR2X1 NOR2_913 (.Y(N2836),.A(N2712),.B(N2769));
NOR2X1 NOR2_914 (.Y(N2837),.A(N2769),.B(N846));
NOR2X1 NOR2_915 (.Y(N2838),.A(N2619),.B(N2769));
NOR2X1 NOR2_916 (.Y(N2841),.A(N2715),.B(N2773));
NOR2X1 NOR2_917 (.Y(N2842),.A(N2773),.B(N894));
NOR2X1 NOR2_918 (.Y(N2843),.A(N2623),.B(N2773));
NOR2X1 NOR2_919 (.Y(N2846),.A(N2718),.B(N2777));
NOR2X1 NOR2_920 (.Y(N2847),.A(N2777),.B(N942));
NOR2X1 NOR2_921 (.Y(N2848),.A(N2627),.B(N2777));
NOR2X1 NOR2_922 (.Y(N2851),.A(N2721),.B(N2781));
NOR2X1 NOR2_923 (.Y(N2852),.A(N2781),.B(N990));
NOR2X1 NOR2_924 (.Y(N2853),.A(N2631),.B(N2781));
NOR2X1 NOR2_925 (.Y(N2856),.A(N2724),.B(N2785));
NOR2X1 NOR2_926 (.Y(N2857),.A(N2785),.B(N1038));
NOR2X1 NOR2_927 (.Y(N2858),.A(N2635),.B(N2785));
NOR2X1 NOR2_928 (.Y(N2861),.A(N2789),.B(N2790));
NOR2X1 NOR2_929 (.Y(N2864),.A(N2794),.B(N2791));
NOR2X1 NOR2_930 (.Y(N2868),.A(N2736),.B(N2797));
NOR2X1 NOR2_931 (.Y(N2869),.A(N2797),.B(N2733));
NOR2X1 NOR2_932 (.Y(N2870),.A(N2801),.B(N2802));
NOR2X1 NOR2_933 (.Y(N2873),.A(N2803),.B(N1233));
NOR2X1 NOR2_934 (.Y(N2877),.A(N2806),.B(N2807));
NOR2X1 NOR2_935 (.Y(N2878),.A(N2811),.B(N2812));
NOR2X1 NOR2_936 (.Y(N2881),.A(N2816),.B(N2817));
NOR2X1 NOR2_937 (.Y(N2884),.A(N2821),.B(N2822));
NOR2X1 NOR2_938 (.Y(N2887),.A(N2826),.B(N2827));
NOR2X1 NOR2_939 (.Y(N2890),.A(N2831),.B(N2832));
NOR2X1 NOR2_940 (.Y(N2893),.A(N2836),.B(N2837));
NOR2X1 NOR2_941 (.Y(N2896),.A(N2841),.B(N2842));
NOR2X1 NOR2_942 (.Y(N2899),.A(N2846),.B(N2847));
NOR2X1 NOR2_943 (.Y(N2902),.A(N2851),.B(N2852));
NOR2X1 NOR2_944 (.Y(N2905),.A(N2856),.B(N2857));
NOR2X1 NOR2_945 (.Y(N2908),.A(N2861),.B(N2858));
NOR2X1 NOR2_946 (.Y(N2912),.A(N2794),.B(N2864));
NOR2X1 NOR2_947 (.Y(N2913),.A(N2864),.B(N2791));
NOR2X1 NOR2_948 (.Y(N2914),.A(N2868),.B(N2869));
NOR2X1 NOR2_949 (.Y(N2917),.A(N2870),.B(N1185));
NOR2X1 NOR2_950 (.Y(N2921),.A(N2803),.B(N2873));
NOR2X1 NOR2_951 (.Y(N2922),.A(N2873),.B(N1233));
NOR2X1 NOR2_952 (.Y(N2923),.A(N2690),.B(N2873));
NOR2X1 NOR2_953 (.Y(N2926),.A(N2878),.B(N2808));
NOR2X1 NOR2_954 (.Y(N2930),.A(N2881),.B(N2813));
NOR2X1 NOR2_955 (.Y(N2934),.A(N2884),.B(N2818));
NOR2X1 NOR2_956 (.Y(N2938),.A(N2887),.B(N2823));
NOR2X1 NOR2_957 (.Y(N2942),.A(N2890),.B(N2828));
NOR2X1 NOR2_958 (.Y(N2946),.A(N2893),.B(N2833));
NOR2X1 NOR2_959 (.Y(N2950),.A(N2896),.B(N2838));
NOR2X1 NOR2_960 (.Y(N2954),.A(N2899),.B(N2843));
NOR2X1 NOR2_961 (.Y(N2958),.A(N2902),.B(N2848));
NOR2X1 NOR2_962 (.Y(N2962),.A(N2905),.B(N2853));
NOR2X1 NOR2_963 (.Y(N2966),.A(N2861),.B(N2908));
NOR2X1 NOR2_964 (.Y(N2967),.A(N2908),.B(N2858));
NOR2X1 NOR2_965 (.Y(N2968),.A(N2912),.B(N2913));
NOR2X1 NOR2_966 (.Y(N2971),.A(N2914),.B(N1137));
NOR2X1 NOR2_967 (.Y(N2975),.A(N2870),.B(N2917));
NOR2X1 NOR2_968 (.Y(N2976),.A(N2917),.B(N1185));
NOR2X1 NOR2_969 (.Y(N2977),.A(N2739),.B(N2917));
NOR2X1 NOR2_970 (.Y(N2980),.A(N2921),.B(N2922));
NOR2X1 NOR2_971 (.Y(N2983),.A(N1281),.B(N2923));
NOR2X1 NOR2_972 (.Y(N2987),.A(N2878),.B(N2926));
NOR2X1 NOR2_973 (.Y(N2988),.A(N2926),.B(N2808));
NOR2X1 NOR2_974 (.Y(N2989),.A(N2881),.B(N2930));
NOR2X1 NOR2_975 (.Y(N2990),.A(N2930),.B(N2813));
NOR2X1 NOR2_976 (.Y(N2991),.A(N2884),.B(N2934));
NOR2X1 NOR2_977 (.Y(N2992),.A(N2934),.B(N2818));
NOR2X1 NOR2_978 (.Y(N2993),.A(N2887),.B(N2938));
NOR2X1 NOR2_979 (.Y(N2994),.A(N2938),.B(N2823));
NOR2X1 NOR2_980 (.Y(N2995),.A(N2890),.B(N2942));
NOR2X1 NOR2_981 (.Y(N2996),.A(N2942),.B(N2828));
NOR2X1 NOR2_982 (.Y(N2997),.A(N2893),.B(N2946));
NOR2X1 NOR2_983 (.Y(N2998),.A(N2946),.B(N2833));
NOR2X1 NOR2_984 (.Y(N2999),.A(N2896),.B(N2950));
NOR2X1 NOR2_985 (.Y(N3000),.A(N2950),.B(N2838));
NOR2X1 NOR2_986 (.Y(N3001),.A(N2899),.B(N2954));
NOR2X1 NOR2_987 (.Y(N3002),.A(N2954),.B(N2843));
NOR2X1 NOR2_988 (.Y(N3003),.A(N2902),.B(N2958));
NOR2X1 NOR2_989 (.Y(N3004),.A(N2958),.B(N2848));
NOR2X1 NOR2_990 (.Y(N3005),.A(N2905),.B(N2962));
NOR2X1 NOR2_991 (.Y(N3006),.A(N2962),.B(N2853));
NOR2X1 NOR2_992 (.Y(N3007),.A(N2966),.B(N2967));
NOR2X1 NOR2_993 (.Y(N3010),.A(N2968),.B(N1089));
NOR2X1 NOR2_994 (.Y(N3014),.A(N2914),.B(N2971));
NOR2X1 NOR2_995 (.Y(N3015),.A(N2971),.B(N1137));
NOR2X1 NOR2_996 (.Y(N3016),.A(N2797),.B(N2971));
NOR2X1 NOR2_997 (.Y(N3019),.A(N2975),.B(N2976));
NOR2X1 NOR2_998 (.Y(N3022),.A(N2980),.B(N2977));
NOR2X1 NOR2_999 (.Y(N3026),.A(N1281),.B(N2983));
NOR2X1 NOR2_1000 (.Y(N3027),.A(N2983),.B(N2923));
NOR2X1 NOR2_1001 (.Y(N3028),.A(N2987),.B(N2988));
NOR2X1 NOR2_1002 (.Y(N3031),.A(N2989),.B(N2990));
NOR2X1 NOR2_1003 (.Y(N3034),.A(N2991),.B(N2992));
NOR2X1 NOR2_1004 (.Y(N3037),.A(N2993),.B(N2994));
NOR2X1 NOR2_1005 (.Y(N3040),.A(N2995),.B(N2996));
NOR2X1 NOR2_1006 (.Y(N3043),.A(N2997),.B(N2998));
NOR2X1 NOR2_1007 (.Y(N3046),.A(N2999),.B(N3000));
NOR2X1 NOR2_1008 (.Y(N3049),.A(N3001),.B(N3002));
NOR2X1 NOR2_1009 (.Y(N3052),.A(N3003),.B(N3004));
NOR2X1 NOR2_1010 (.Y(N3055),.A(N3005),.B(N3006));
NOR2X1 NOR2_1011 (.Y(N3058),.A(N3007),.B(N1041));
NOR2X1 NOR2_1012 (.Y(N3062),.A(N2968),.B(N3010));
NOR2X1 NOR2_1013 (.Y(N3063),.A(N3010),.B(N1089));
NOR2X1 NOR2_1014 (.Y(N3064),.A(N2864),.B(N3010));
NOR2X1 NOR2_1015 (.Y(N3067),.A(N3014),.B(N3015));
NOR2X1 NOR2_1016 (.Y(N3070),.A(N3019),.B(N3016));
NOR2X1 NOR2_1017 (.Y(N3074),.A(N2980),.B(N3022));
NOR2X1 NOR2_1018 (.Y(N3075),.A(N3022),.B(N2977));
NOR2X1 NOR2_1019 (.Y(N3076),.A(N3026),.B(N3027));
NOR2X1 NOR2_1020 (.Y(N3079),.A(N3028),.B(N561));
NOR2X1 NOR2_1021 (.Y(N3083),.A(N3031),.B(N609));
NOR2X1 NOR2_1022 (.Y(N3087),.A(N3034),.B(N657));
NOR2X1 NOR2_1023 (.Y(N3091),.A(N3037),.B(N705));
NOR2X1 NOR2_1024 (.Y(N3095),.A(N3040),.B(N753));
NOR2X1 NOR2_1025 (.Y(N3099),.A(N3043),.B(N801));
NOR2X1 NOR2_1026 (.Y(N3103),.A(N3046),.B(N849));
NOR2X1 NOR2_1027 (.Y(N3107),.A(N3049),.B(N897));
NOR2X1 NOR2_1028 (.Y(N3111),.A(N3052),.B(N945));
NOR2X1 NOR2_1029 (.Y(N3115),.A(N3055),.B(N993));
NOR2X1 NOR2_1030 (.Y(N3119),.A(N3007),.B(N3058));
NOR2X1 NOR2_1031 (.Y(N3120),.A(N3058),.B(N1041));
NOR2X1 NOR2_1032 (.Y(N3121),.A(N2908),.B(N3058));
NOR2X1 NOR2_1033 (.Y(N3124),.A(N3062),.B(N3063));
NOR2X1 NOR2_1034 (.Y(N3127),.A(N3067),.B(N3064));
NOR2X1 NOR2_1035 (.Y(N3131),.A(N3019),.B(N3070));
NOR2X1 NOR2_1036 (.Y(N3132),.A(N3070),.B(N3016));
NOR2X1 NOR2_1037 (.Y(N3133),.A(N3074),.B(N3075));
NOR2X1 NOR2_1038 (.Y(N3136),.A(N3076),.B(N1236));
NOR2X1 NOR2_1039 (.Y(N3140),.A(N3028),.B(N3079));
NOR2X1 NOR2_1040 (.Y(N3141),.A(N3079),.B(N561));
NOR2X1 NOR2_1041 (.Y(N3142),.A(N2926),.B(N3079));
NOR2X1 NOR2_1042 (.Y(N3145),.A(N3031),.B(N3083));
NOR2X1 NOR2_1043 (.Y(N3146),.A(N3083),.B(N609));
NOR2X1 NOR2_1044 (.Y(N3147),.A(N2930),.B(N3083));
NOR2X1 NOR2_1045 (.Y(N3150),.A(N3034),.B(N3087));
NOR2X1 NOR2_1046 (.Y(N3151),.A(N3087),.B(N657));
NOR2X1 NOR2_1047 (.Y(N3152),.A(N2934),.B(N3087));
NOR2X1 NOR2_1048 (.Y(N3155),.A(N3037),.B(N3091));
NOR2X1 NOR2_1049 (.Y(N3156),.A(N3091),.B(N705));
NOR2X1 NOR2_1050 (.Y(N3157),.A(N2938),.B(N3091));
NOR2X1 NOR2_1051 (.Y(N3160),.A(N3040),.B(N3095));
NOR2X1 NOR2_1052 (.Y(N3161),.A(N3095),.B(N753));
NOR2X1 NOR2_1053 (.Y(N3162),.A(N2942),.B(N3095));
NOR2X1 NOR2_1054 (.Y(N3165),.A(N3043),.B(N3099));
NOR2X1 NOR2_1055 (.Y(N3166),.A(N3099),.B(N801));
NOR2X1 NOR2_1056 (.Y(N3167),.A(N2946),.B(N3099));
NOR2X1 NOR2_1057 (.Y(N3170),.A(N3046),.B(N3103));
NOR2X1 NOR2_1058 (.Y(N3171),.A(N3103),.B(N849));
NOR2X1 NOR2_1059 (.Y(N3172),.A(N2950),.B(N3103));
NOR2X1 NOR2_1060 (.Y(N3175),.A(N3049),.B(N3107));
NOR2X1 NOR2_1061 (.Y(N3176),.A(N3107),.B(N897));
NOR2X1 NOR2_1062 (.Y(N3177),.A(N2954),.B(N3107));
NOR2X1 NOR2_1063 (.Y(N3180),.A(N3052),.B(N3111));
NOR2X1 NOR2_1064 (.Y(N3181),.A(N3111),.B(N945));
NOR2X1 NOR2_1065 (.Y(N3182),.A(N2958),.B(N3111));
NOR2X1 NOR2_1066 (.Y(N3185),.A(N3055),.B(N3115));
NOR2X1 NOR2_1067 (.Y(N3186),.A(N3115),.B(N993));
NOR2X1 NOR2_1068 (.Y(N3187),.A(N2962),.B(N3115));
NOR2X1 NOR2_1069 (.Y(N3190),.A(N3119),.B(N3120));
NOR2X1 NOR2_1070 (.Y(N3193),.A(N3124),.B(N3121));
NOR2X1 NOR2_1071 (.Y(N3197),.A(N3067),.B(N3127));
NOR2X1 NOR2_1072 (.Y(N3198),.A(N3127),.B(N3064));
NOR2X1 NOR2_1073 (.Y(N3199),.A(N3131),.B(N3132));
NOR2X1 NOR2_1074 (.Y(N3202),.A(N3133),.B(N1188));
NOR2X1 NOR2_1075 (.Y(N3206),.A(N3076),.B(N3136));
NOR2X1 NOR2_1076 (.Y(N3207),.A(N3136),.B(N1236));
NOR2X1 NOR2_1077 (.Y(N3208),.A(N2983),.B(N3136));
NOR2X1 NOR2_1078 (.Y(N3211),.A(N3140),.B(N3141));
NOR2X1 NOR2_1079 (.Y(N3212),.A(N3145),.B(N3146));
NOR2X1 NOR2_1080 (.Y(N3215),.A(N3150),.B(N3151));
NOR2X1 NOR2_1081 (.Y(N3218),.A(N3155),.B(N3156));
NOR2X1 NOR2_1082 (.Y(N3221),.A(N3160),.B(N3161));
NOR2X1 NOR2_1083 (.Y(N3224),.A(N3165),.B(N3166));
NOR2X1 NOR2_1084 (.Y(N3227),.A(N3170),.B(N3171));
NOR2X1 NOR2_1085 (.Y(N3230),.A(N3175),.B(N3176));
NOR2X1 NOR2_1086 (.Y(N3233),.A(N3180),.B(N3181));
NOR2X1 NOR2_1087 (.Y(N3236),.A(N3185),.B(N3186));
NOR2X1 NOR2_1088 (.Y(N3239),.A(N3190),.B(N3187));
NOR2X1 NOR2_1089 (.Y(N3243),.A(N3124),.B(N3193));
NOR2X1 NOR2_1090 (.Y(N3244),.A(N3193),.B(N3121));
NOR2X1 NOR2_1091 (.Y(N3245),.A(N3197),.B(N3198));
NOR2X1 NOR2_1092 (.Y(N3248),.A(N3199),.B(N1140));
NOR2X1 NOR2_1093 (.Y(N3252),.A(N3133),.B(N3202));
NOR2X1 NOR2_1094 (.Y(N3253),.A(N3202),.B(N1188));
NOR2X1 NOR2_1095 (.Y(N3254),.A(N3022),.B(N3202));
NOR2X1 NOR2_1096 (.Y(N3257),.A(N3206),.B(N3207));
NOR2X1 NOR2_1097 (.Y(N3260),.A(N1284),.B(N3208));
NOR2X1 NOR2_1098 (.Y(N3264),.A(N3212),.B(N3142));
NOR2X1 NOR2_1099 (.Y(N3268),.A(N3215),.B(N3147));
NOR2X1 NOR2_1100 (.Y(N3272),.A(N3218),.B(N3152));
NOR2X1 NOR2_1101 (.Y(N3276),.A(N3221),.B(N3157));
NOR2X1 NOR2_1102 (.Y(N3280),.A(N3224),.B(N3162));
NOR2X1 NOR2_1103 (.Y(N3284),.A(N3227),.B(N3167));
NOR2X1 NOR2_1104 (.Y(N3288),.A(N3230),.B(N3172));
NOR2X1 NOR2_1105 (.Y(N3292),.A(N3233),.B(N3177));
NOR2X1 NOR2_1106 (.Y(N3296),.A(N3236),.B(N3182));
NOR2X1 NOR2_1107 (.Y(N3300),.A(N3190),.B(N3239));
NOR2X1 NOR2_1108 (.Y(N3301),.A(N3239),.B(N3187));
NOR2X1 NOR2_1109 (.Y(N3302),.A(N3243),.B(N3244));
NOR2X1 NOR2_1110 (.Y(N3305),.A(N3245),.B(N1092));
NOR2X1 NOR2_1111 (.Y(N3309),.A(N3199),.B(N3248));
NOR2X1 NOR2_1112 (.Y(N3310),.A(N3248),.B(N1140));
NOR2X1 NOR2_1113 (.Y(N3311),.A(N3070),.B(N3248));
NOR2X1 NOR2_1114 (.Y(N3314),.A(N3252),.B(N3253));
NOR2X1 NOR2_1115 (.Y(N3317),.A(N3257),.B(N3254));
NOR2X1 NOR2_1116 (.Y(N3321),.A(N1284),.B(N3260));
NOR2X1 NOR2_1117 (.Y(N3322),.A(N3260),.B(N3208));
NOR2X1 NOR2_1118 (.Y(N3323),.A(N3212),.B(N3264));
NOR2X1 NOR2_1119 (.Y(N3324),.A(N3264),.B(N3142));
NOR2X1 NOR2_1120 (.Y(N3325),.A(N3215),.B(N3268));
NOR2X1 NOR2_1121 (.Y(N3326),.A(N3268),.B(N3147));
NOR2X1 NOR2_1122 (.Y(N3327),.A(N3218),.B(N3272));
NOR2X1 NOR2_1123 (.Y(N3328),.A(N3272),.B(N3152));
NOR2X1 NOR2_1124 (.Y(N3329),.A(N3221),.B(N3276));
NOR2X1 NOR2_1125 (.Y(N3330),.A(N3276),.B(N3157));
NOR2X1 NOR2_1126 (.Y(N3331),.A(N3224),.B(N3280));
NOR2X1 NOR2_1127 (.Y(N3332),.A(N3280),.B(N3162));
NOR2X1 NOR2_1128 (.Y(N3333),.A(N3227),.B(N3284));
NOR2X1 NOR2_1129 (.Y(N3334),.A(N3284),.B(N3167));
NOR2X1 NOR2_1130 (.Y(N3335),.A(N3230),.B(N3288));
NOR2X1 NOR2_1131 (.Y(N3336),.A(N3288),.B(N3172));
NOR2X1 NOR2_1132 (.Y(N3337),.A(N3233),.B(N3292));
NOR2X1 NOR2_1133 (.Y(N3338),.A(N3292),.B(N3177));
NOR2X1 NOR2_1134 (.Y(N3339),.A(N3236),.B(N3296));
NOR2X1 NOR2_1135 (.Y(N3340),.A(N3296),.B(N3182));
NOR2X1 NOR2_1136 (.Y(N3341),.A(N3300),.B(N3301));
NOR2X1 NOR2_1137 (.Y(N3344),.A(N3302),.B(N1044));
NOR2X1 NOR2_1138 (.Y(N3348),.A(N3245),.B(N3305));
NOR2X1 NOR2_1139 (.Y(N3349),.A(N3305),.B(N1092));
NOR2X1 NOR2_1140 (.Y(N3350),.A(N3127),.B(N3305));
NOR2X1 NOR2_1141 (.Y(N3353),.A(N3309),.B(N3310));
NOR2X1 NOR2_1142 (.Y(N3356),.A(N3314),.B(N3311));
NOR2X1 NOR2_1143 (.Y(N3360),.A(N3257),.B(N3317));
NOR2X1 NOR2_1144 (.Y(N3361),.A(N3317),.B(N3254));
NOR2X1 NOR2_1145 (.Y(N3362),.A(N3321),.B(N3322));
NOR2X1 NOR2_1146 (.Y(N3365),.A(N3323),.B(N3324));
NOR2X1 NOR2_1147 (.Y(N3368),.A(N3325),.B(N3326));
NOR2X1 NOR2_1148 (.Y(N3371),.A(N3327),.B(N3328));
NOR2X1 NOR2_1149 (.Y(N3374),.A(N3329),.B(N3330));
NOR2X1 NOR2_1150 (.Y(N3377),.A(N3331),.B(N3332));
NOR2X1 NOR2_1151 (.Y(N3380),.A(N3333),.B(N3334));
NOR2X1 NOR2_1152 (.Y(N3383),.A(N3335),.B(N3336));
NOR2X1 NOR2_1153 (.Y(N3386),.A(N3337),.B(N3338));
NOR2X1 NOR2_1154 (.Y(N3389),.A(N3339),.B(N3340));
NOR2X1 NOR2_1155 (.Y(N3392),.A(N3341),.B(N996));
NOR2X1 NOR2_1156 (.Y(N3396),.A(N3302),.B(N3344));
NOR2X1 NOR2_1157 (.Y(N3397),.A(N3344),.B(N1044));
NOR2X1 NOR2_1158 (.Y(N3398),.A(N3193),.B(N3344));
NOR2X1 NOR2_1159 (.Y(N3401),.A(N3348),.B(N3349));
NOR2X1 NOR2_1160 (.Y(N3404),.A(N3353),.B(N3350));
NOR2X1 NOR2_1161 (.Y(N3408),.A(N3314),.B(N3356));
NOR2X1 NOR2_1162 (.Y(N3409),.A(N3356),.B(N3311));
NOR2X1 NOR2_1163 (.Y(N3410),.A(N3360),.B(N3361));
NOR2X1 NOR2_1164 (.Y(N3413),.A(N3362),.B(N1239));
NOR2X1 NOR2_1165 (.Y(N3417),.A(N3365),.B(N564));
NOR2X1 NOR2_1166 (.Y(N3421),.A(N3368),.B(N612));
NOR2X1 NOR2_1167 (.Y(N3425),.A(N3371),.B(N660));
NOR2X1 NOR2_1168 (.Y(N3429),.A(N3374),.B(N708));
NOR2X1 NOR2_1169 (.Y(N3433),.A(N3377),.B(N756));
NOR2X1 NOR2_1170 (.Y(N3437),.A(N3380),.B(N804));
NOR2X1 NOR2_1171 (.Y(N3441),.A(N3383),.B(N852));
NOR2X1 NOR2_1172 (.Y(N3445),.A(N3386),.B(N900));
NOR2X1 NOR2_1173 (.Y(N3449),.A(N3389),.B(N948));
NOR2X1 NOR2_1174 (.Y(N3453),.A(N3341),.B(N3392));
NOR2X1 NOR2_1175 (.Y(N3454),.A(N3392),.B(N996));
NOR2X1 NOR2_1176 (.Y(N3455),.A(N3239),.B(N3392));
NOR2X1 NOR2_1177 (.Y(N3458),.A(N3396),.B(N3397));
NOR2X1 NOR2_1178 (.Y(N3461),.A(N3401),.B(N3398));
NOR2X1 NOR2_1179 (.Y(N3465),.A(N3353),.B(N3404));
NOR2X1 NOR2_1180 (.Y(N3466),.A(N3404),.B(N3350));
NOR2X1 NOR2_1181 (.Y(N3467),.A(N3408),.B(N3409));
NOR2X1 NOR2_1182 (.Y(N3470),.A(N3410),.B(N1191));
NOR2X1 NOR2_1183 (.Y(N3474),.A(N3362),.B(N3413));
NOR2X1 NOR2_1184 (.Y(N3475),.A(N3413),.B(N1239));
NOR2X1 NOR2_1185 (.Y(N3476),.A(N3260),.B(N3413));
NOR2X1 NOR2_1186 (.Y(N3479),.A(N3365),.B(N3417));
NOR2X1 NOR2_1187 (.Y(N3480),.A(N3417),.B(N564));
NOR2X1 NOR2_1188 (.Y(N3481),.A(N3264),.B(N3417));
NOR2X1 NOR2_1189 (.Y(N3484),.A(N3368),.B(N3421));
NOR2X1 NOR2_1190 (.Y(N3485),.A(N3421),.B(N612));
NOR2X1 NOR2_1191 (.Y(N3486),.A(N3268),.B(N3421));
NOR2X1 NOR2_1192 (.Y(N3489),.A(N3371),.B(N3425));
NOR2X1 NOR2_1193 (.Y(N3490),.A(N3425),.B(N660));
NOR2X1 NOR2_1194 (.Y(N3491),.A(N3272),.B(N3425));
NOR2X1 NOR2_1195 (.Y(N3494),.A(N3374),.B(N3429));
NOR2X1 NOR2_1196 (.Y(N3495),.A(N3429),.B(N708));
NOR2X1 NOR2_1197 (.Y(N3496),.A(N3276),.B(N3429));
NOR2X1 NOR2_1198 (.Y(N3499),.A(N3377),.B(N3433));
NOR2X1 NOR2_1199 (.Y(N3500),.A(N3433),.B(N756));
NOR2X1 NOR2_1200 (.Y(N3501),.A(N3280),.B(N3433));
NOR2X1 NOR2_1201 (.Y(N3504),.A(N3380),.B(N3437));
NOR2X1 NOR2_1202 (.Y(N3505),.A(N3437),.B(N804));
NOR2X1 NOR2_1203 (.Y(N3506),.A(N3284),.B(N3437));
NOR2X1 NOR2_1204 (.Y(N3509),.A(N3383),.B(N3441));
NOR2X1 NOR2_1205 (.Y(N3510),.A(N3441),.B(N852));
NOR2X1 NOR2_1206 (.Y(N3511),.A(N3288),.B(N3441));
NOR2X1 NOR2_1207 (.Y(N3514),.A(N3386),.B(N3445));
NOR2X1 NOR2_1208 (.Y(N3515),.A(N3445),.B(N900));
NOR2X1 NOR2_1209 (.Y(N3516),.A(N3292),.B(N3445));
NOR2X1 NOR2_1210 (.Y(N3519),.A(N3389),.B(N3449));
NOR2X1 NOR2_1211 (.Y(N3520),.A(N3449),.B(N948));
NOR2X1 NOR2_1212 (.Y(N3521),.A(N3296),.B(N3449));
NOR2X1 NOR2_1213 (.Y(N3524),.A(N3453),.B(N3454));
NOR2X1 NOR2_1214 (.Y(N3527),.A(N3458),.B(N3455));
NOR2X1 NOR2_1215 (.Y(N3531),.A(N3401),.B(N3461));
NOR2X1 NOR2_1216 (.Y(N3532),.A(N3461),.B(N3398));
NOR2X1 NOR2_1217 (.Y(N3533),.A(N3465),.B(N3466));
NOR2X1 NOR2_1218 (.Y(N3536),.A(N3467),.B(N1143));
NOR2X1 NOR2_1219 (.Y(N3540),.A(N3410),.B(N3470));
NOR2X1 NOR2_1220 (.Y(N3541),.A(N3470),.B(N1191));
NOR2X1 NOR2_1221 (.Y(N3542),.A(N3317),.B(N3470));
NOR2X1 NOR2_1222 (.Y(N3545),.A(N3474),.B(N3475));
NOR2X1 NOR2_1223 (.Y(N3548),.A(N1287),.B(N3476));
NOR2X1 NOR2_1224 (.Y(N3552),.A(N3479),.B(N3480));
NOR2X1 NOR2_1225 (.Y(N3553),.A(N3484),.B(N3485));
NOR2X1 NOR2_1226 (.Y(N3556),.A(N3489),.B(N3490));
NOR2X1 NOR2_1227 (.Y(N3559),.A(N3494),.B(N3495));
NOR2X1 NOR2_1228 (.Y(N3562),.A(N3499),.B(N3500));
NOR2X1 NOR2_1229 (.Y(N3565),.A(N3504),.B(N3505));
NOR2X1 NOR2_1230 (.Y(N3568),.A(N3509),.B(N3510));
NOR2X1 NOR2_1231 (.Y(N3571),.A(N3514),.B(N3515));
NOR2X1 NOR2_1232 (.Y(N3574),.A(N3519),.B(N3520));
NOR2X1 NOR2_1233 (.Y(N3577),.A(N3524),.B(N3521));
NOR2X1 NOR2_1234 (.Y(N3581),.A(N3458),.B(N3527));
NOR2X1 NOR2_1235 (.Y(N3582),.A(N3527),.B(N3455));
NOR2X1 NOR2_1236 (.Y(N3583),.A(N3531),.B(N3532));
NOR2X1 NOR2_1237 (.Y(N3586),.A(N3533),.B(N1095));
NOR2X1 NOR2_1238 (.Y(N3590),.A(N3467),.B(N3536));
NOR2X1 NOR2_1239 (.Y(N3591),.A(N3536),.B(N1143));
NOR2X1 NOR2_1240 (.Y(N3592),.A(N3356),.B(N3536));
NOR2X1 NOR2_1241 (.Y(N3595),.A(N3540),.B(N3541));
NOR2X1 NOR2_1242 (.Y(N3598),.A(N3545),.B(N3542));
NOR2X1 NOR2_1243 (.Y(N3602),.A(N1287),.B(N3548));
NOR2X1 NOR2_1244 (.Y(N3603),.A(N3548),.B(N3476));
NOR2X1 NOR2_1245 (.Y(N3604),.A(N3553),.B(N3481));
NOR2X1 NOR2_1246 (.Y(N3608),.A(N3556),.B(N3486));
NOR2X1 NOR2_1247 (.Y(N3612),.A(N3559),.B(N3491));
NOR2X1 NOR2_1248 (.Y(N3616),.A(N3562),.B(N3496));
NOR2X1 NOR2_1249 (.Y(N3620),.A(N3565),.B(N3501));
NOR2X1 NOR2_1250 (.Y(N3624),.A(N3568),.B(N3506));
NOR2X1 NOR2_1251 (.Y(N3628),.A(N3571),.B(N3511));
NOR2X1 NOR2_1252 (.Y(N3632),.A(N3574),.B(N3516));
NOR2X1 NOR2_1253 (.Y(N3636),.A(N3524),.B(N3577));
NOR2X1 NOR2_1254 (.Y(N3637),.A(N3577),.B(N3521));
NOR2X1 NOR2_1255 (.Y(N3638),.A(N3581),.B(N3582));
NOR2X1 NOR2_1256 (.Y(N3641),.A(N3583),.B(N1047));
NOR2X1 NOR2_1257 (.Y(N3645),.A(N3533),.B(N3586));
NOR2X1 NOR2_1258 (.Y(N3646),.A(N3586),.B(N1095));
NOR2X1 NOR2_1259 (.Y(N3647),.A(N3404),.B(N3586));
NOR2X1 NOR2_1260 (.Y(N3650),.A(N3590),.B(N3591));
NOR2X1 NOR2_1261 (.Y(N3653),.A(N3595),.B(N3592));
NOR2X1 NOR2_1262 (.Y(N3657),.A(N3545),.B(N3598));
NOR2X1 NOR2_1263 (.Y(N3658),.A(N3598),.B(N3542));
NOR2X1 NOR2_1264 (.Y(N3659),.A(N3602),.B(N3603));
NOR2X1 NOR2_1265 (.Y(N3662),.A(N3553),.B(N3604));
NOR2X1 NOR2_1266 (.Y(N3663),.A(N3604),.B(N3481));
NOR2X1 NOR2_1267 (.Y(N3664),.A(N3556),.B(N3608));
NOR2X1 NOR2_1268 (.Y(N3665),.A(N3608),.B(N3486));
NOR2X1 NOR2_1269 (.Y(N3666),.A(N3559),.B(N3612));
NOR2X1 NOR2_1270 (.Y(N3667),.A(N3612),.B(N3491));
NOR2X1 NOR2_1271 (.Y(N3668),.A(N3562),.B(N3616));
NOR2X1 NOR2_1272 (.Y(N3669),.A(N3616),.B(N3496));
NOR2X1 NOR2_1273 (.Y(N3670),.A(N3565),.B(N3620));
NOR2X1 NOR2_1274 (.Y(N3671),.A(N3620),.B(N3501));
NOR2X1 NOR2_1275 (.Y(N3672),.A(N3568),.B(N3624));
NOR2X1 NOR2_1276 (.Y(N3673),.A(N3624),.B(N3506));
NOR2X1 NOR2_1277 (.Y(N3674),.A(N3571),.B(N3628));
NOR2X1 NOR2_1278 (.Y(N3675),.A(N3628),.B(N3511));
NOR2X1 NOR2_1279 (.Y(N3676),.A(N3574),.B(N3632));
NOR2X1 NOR2_1280 (.Y(N3677),.A(N3632),.B(N3516));
NOR2X1 NOR2_1281 (.Y(N3678),.A(N3636),.B(N3637));
NOR2X1 NOR2_1282 (.Y(N3681),.A(N3638),.B(N999));
NOR2X1 NOR2_1283 (.Y(N3685),.A(N3583),.B(N3641));
NOR2X1 NOR2_1284 (.Y(N3686),.A(N3641),.B(N1047));
NOR2X1 NOR2_1285 (.Y(N3687),.A(N3461),.B(N3641));
NOR2X1 NOR2_1286 (.Y(N3690),.A(N3645),.B(N3646));
NOR2X1 NOR2_1287 (.Y(N3693),.A(N3650),.B(N3647));
NOR2X1 NOR2_1288 (.Y(N3697),.A(N3595),.B(N3653));
NOR2X1 NOR2_1289 (.Y(N3698),.A(N3653),.B(N3592));
NOR2X1 NOR2_1290 (.Y(N3699),.A(N3657),.B(N3658));
NOR2X1 NOR2_1291 (.Y(N3702),.A(N3659),.B(N1242));
NOR2X1 NOR2_1292 (.Y(N3706),.A(N3662),.B(N3663));
NOR2X1 NOR2_1293 (.Y(N3709),.A(N3664),.B(N3665));
NOR2X1 NOR2_1294 (.Y(N3712),.A(N3666),.B(N3667));
NOR2X1 NOR2_1295 (.Y(N3715),.A(N3668),.B(N3669));
NOR2X1 NOR2_1296 (.Y(N3718),.A(N3670),.B(N3671));
NOR2X1 NOR2_1297 (.Y(N3721),.A(N3672),.B(N3673));
NOR2X1 NOR2_1298 (.Y(N3724),.A(N3674),.B(N3675));
NOR2X1 NOR2_1299 (.Y(N3727),.A(N3676),.B(N3677));
NOR2X1 NOR2_1300 (.Y(N3730),.A(N3678),.B(N951));
NOR2X1 NOR2_1301 (.Y(N3734),.A(N3638),.B(N3681));
NOR2X1 NOR2_1302 (.Y(N3735),.A(N3681),.B(N999));
NOR2X1 NOR2_1303 (.Y(N3736),.A(N3527),.B(N3681));
NOR2X1 NOR2_1304 (.Y(N3739),.A(N3685),.B(N3686));
NOR2X1 NOR2_1305 (.Y(N3742),.A(N3690),.B(N3687));
NOR2X1 NOR2_1306 (.Y(N3746),.A(N3650),.B(N3693));
NOR2X1 NOR2_1307 (.Y(N3747),.A(N3693),.B(N3647));
NOR2X1 NOR2_1308 (.Y(N3748),.A(N3697),.B(N3698));
NOR2X1 NOR2_1309 (.Y(N3751),.A(N3699),.B(N1194));
NOR2X1 NOR2_1310 (.Y(N3755),.A(N3659),.B(N3702));
NOR2X1 NOR2_1311 (.Y(N3756),.A(N3702),.B(N1242));
NOR2X1 NOR2_1312 (.Y(N3757),.A(N3548),.B(N3702));
NOR2X1 NOR2_1313 (.Y(N3760),.A(N3706),.B(N567));
NOR2X1 NOR2_1314 (.Y(N3764),.A(N3709),.B(N615));
NOR2X1 NOR2_1315 (.Y(N3768),.A(N3712),.B(N663));
NOR2X1 NOR2_1316 (.Y(N3772),.A(N3715),.B(N711));
NOR2X1 NOR2_1317 (.Y(N3776),.A(N3718),.B(N759));
NOR2X1 NOR2_1318 (.Y(N3780),.A(N3721),.B(N807));
NOR2X1 NOR2_1319 (.Y(N3784),.A(N3724),.B(N855));
NOR2X1 NOR2_1320 (.Y(N3788),.A(N3727),.B(N903));
NOR2X1 NOR2_1321 (.Y(N3792),.A(N3678),.B(N3730));
NOR2X1 NOR2_1322 (.Y(N3793),.A(N3730),.B(N951));
NOR2X1 NOR2_1323 (.Y(N3794),.A(N3577),.B(N3730));
NOR2X1 NOR2_1324 (.Y(N3797),.A(N3734),.B(N3735));
NOR2X1 NOR2_1325 (.Y(N3800),.A(N3739),.B(N3736));
NOR2X1 NOR2_1326 (.Y(N3804),.A(N3690),.B(N3742));
NOR2X1 NOR2_1327 (.Y(N3805),.A(N3742),.B(N3687));
NOR2X1 NOR2_1328 (.Y(N3806),.A(N3746),.B(N3747));
NOR2X1 NOR2_1329 (.Y(N3809),.A(N3748),.B(N1146));
NOR2X1 NOR2_1330 (.Y(N3813),.A(N3699),.B(N3751));
NOR2X1 NOR2_1331 (.Y(N3814),.A(N3751),.B(N1194));
NOR2X1 NOR2_1332 (.Y(N3815),.A(N3598),.B(N3751));
NOR2X1 NOR2_1333 (.Y(N3818),.A(N3755),.B(N3756));
NOR2X1 NOR2_1334 (.Y(N3821),.A(N1290),.B(N3757));
NOR2X1 NOR2_1335 (.Y(N3825),.A(N3706),.B(N3760));
NOR2X1 NOR2_1336 (.Y(N3826),.A(N3760),.B(N567));
NOR2X1 NOR2_1337 (.Y(N3827),.A(N3604),.B(N3760));
NOR2X1 NOR2_1338 (.Y(N3830),.A(N3709),.B(N3764));
NOR2X1 NOR2_1339 (.Y(N3831),.A(N3764),.B(N615));
NOR2X1 NOR2_1340 (.Y(N3832),.A(N3608),.B(N3764));
NOR2X1 NOR2_1341 (.Y(N3835),.A(N3712),.B(N3768));
NOR2X1 NOR2_1342 (.Y(N3836),.A(N3768),.B(N663));
NOR2X1 NOR2_1343 (.Y(N3837),.A(N3612),.B(N3768));
NOR2X1 NOR2_1344 (.Y(N3840),.A(N3715),.B(N3772));
NOR2X1 NOR2_1345 (.Y(N3841),.A(N3772),.B(N711));
NOR2X1 NOR2_1346 (.Y(N3842),.A(N3616),.B(N3772));
NOR2X1 NOR2_1347 (.Y(N3845),.A(N3718),.B(N3776));
NOR2X1 NOR2_1348 (.Y(N3846),.A(N3776),.B(N759));
NOR2X1 NOR2_1349 (.Y(N3847),.A(N3620),.B(N3776));
NOR2X1 NOR2_1350 (.Y(N3850),.A(N3721),.B(N3780));
NOR2X1 NOR2_1351 (.Y(N3851),.A(N3780),.B(N807));
NOR2X1 NOR2_1352 (.Y(N3852),.A(N3624),.B(N3780));
NOR2X1 NOR2_1353 (.Y(N3855),.A(N3724),.B(N3784));
NOR2X1 NOR2_1354 (.Y(N3856),.A(N3784),.B(N855));
NOR2X1 NOR2_1355 (.Y(N3857),.A(N3628),.B(N3784));
NOR2X1 NOR2_1356 (.Y(N3860),.A(N3727),.B(N3788));
NOR2X1 NOR2_1357 (.Y(N3861),.A(N3788),.B(N903));
NOR2X1 NOR2_1358 (.Y(N3862),.A(N3632),.B(N3788));
NOR2X1 NOR2_1359 (.Y(N3865),.A(N3792),.B(N3793));
NOR2X1 NOR2_1360 (.Y(N3868),.A(N3797),.B(N3794));
NOR2X1 NOR2_1361 (.Y(N3872),.A(N3739),.B(N3800));
NOR2X1 NOR2_1362 (.Y(N3873),.A(N3800),.B(N3736));
NOR2X1 NOR2_1363 (.Y(N3874),.A(N3804),.B(N3805));
NOR2X1 NOR2_1364 (.Y(N3877),.A(N3806),.B(N1098));
NOR2X1 NOR2_1365 (.Y(N3881),.A(N3748),.B(N3809));
NOR2X1 NOR2_1366 (.Y(N3882),.A(N3809),.B(N1146));
NOR2X1 NOR2_1367 (.Y(N3883),.A(N3653),.B(N3809));
NOR2X1 NOR2_1368 (.Y(N3886),.A(N3813),.B(N3814));
NOR2X1 NOR2_1369 (.Y(N3889),.A(N3818),.B(N3815));
NOR2X1 NOR2_1370 (.Y(N3893),.A(N1290),.B(N3821));
NOR2X1 NOR2_1371 (.Y(N3894),.A(N3821),.B(N3757));
NOR2X1 NOR2_1372 (.Y(N3895),.A(N3825),.B(N3826));
NOR2X1 NOR2_1373 (.Y(N3896),.A(N3830),.B(N3831));
NOR2X1 NOR2_1374 (.Y(N3899),.A(N3835),.B(N3836));
NOR2X1 NOR2_1375 (.Y(N3902),.A(N3840),.B(N3841));
NOR2X1 NOR2_1376 (.Y(N3905),.A(N3845),.B(N3846));
NOR2X1 NOR2_1377 (.Y(N3908),.A(N3850),.B(N3851));
NOR2X1 NOR2_1378 (.Y(N3911),.A(N3855),.B(N3856));
NOR2X1 NOR2_1379 (.Y(N3914),.A(N3860),.B(N3861));
NOR2X1 NOR2_1380 (.Y(N3917),.A(N3865),.B(N3862));
NOR2X1 NOR2_1381 (.Y(N3921),.A(N3797),.B(N3868));
NOR2X1 NOR2_1382 (.Y(N3922),.A(N3868),.B(N3794));
NOR2X1 NOR2_1383 (.Y(N3923),.A(N3872),.B(N3873));
NOR2X1 NOR2_1384 (.Y(N3926),.A(N3874),.B(N1050));
NOR2X1 NOR2_1385 (.Y(N3930),.A(N3806),.B(N3877));
NOR2X1 NOR2_1386 (.Y(N3931),.A(N3877),.B(N1098));
NOR2X1 NOR2_1387 (.Y(N3932),.A(N3693),.B(N3877));
NOR2X1 NOR2_1388 (.Y(N3935),.A(N3881),.B(N3882));
NOR2X1 NOR2_1389 (.Y(N3938),.A(N3886),.B(N3883));
NOR2X1 NOR2_1390 (.Y(N3942),.A(N3818),.B(N3889));
NOR2X1 NOR2_1391 (.Y(N3943),.A(N3889),.B(N3815));
NOR2X1 NOR2_1392 (.Y(N3944),.A(N3893),.B(N3894));
NOR2X1 NOR2_1393 (.Y(N3947),.A(N3896),.B(N3827));
NOR2X1 NOR2_1394 (.Y(N3951),.A(N3899),.B(N3832));
NOR2X1 NOR2_1395 (.Y(N3955),.A(N3902),.B(N3837));
NOR2X1 NOR2_1396 (.Y(N3959),.A(N3905),.B(N3842));
NOR2X1 NOR2_1397 (.Y(N3963),.A(N3908),.B(N3847));
NOR2X1 NOR2_1398 (.Y(N3967),.A(N3911),.B(N3852));
NOR2X1 NOR2_1399 (.Y(N3971),.A(N3914),.B(N3857));
NOR2X1 NOR2_1400 (.Y(N3975),.A(N3865),.B(N3917));
NOR2X1 NOR2_1401 (.Y(N3976),.A(N3917),.B(N3862));
NOR2X1 NOR2_1402 (.Y(N3977),.A(N3921),.B(N3922));
NOR2X1 NOR2_1403 (.Y(N3980),.A(N3923),.B(N1002));
NOR2X1 NOR2_1404 (.Y(N3984),.A(N3874),.B(N3926));
NOR2X1 NOR2_1405 (.Y(N3985),.A(N3926),.B(N1050));
NOR2X1 NOR2_1406 (.Y(N3986),.A(N3742),.B(N3926));
NOR2X1 NOR2_1407 (.Y(N3989),.A(N3930),.B(N3931));
NOR2X1 NOR2_1408 (.Y(N3992),.A(N3935),.B(N3932));
NOR2X1 NOR2_1409 (.Y(N3996),.A(N3886),.B(N3938));
NOR2X1 NOR2_1410 (.Y(N3997),.A(N3938),.B(N3883));
NOR2X1 NOR2_1411 (.Y(N3998),.A(N3942),.B(N3943));
NOR2X1 NOR2_1412 (.Y(N4001),.A(N3944),.B(N1245));
NOR2X1 NOR2_1413 (.Y(N4005),.A(N3896),.B(N3947));
NOR2X1 NOR2_1414 (.Y(N4006),.A(N3947),.B(N3827));
NOR2X1 NOR2_1415 (.Y(N4007),.A(N3899),.B(N3951));
NOR2X1 NOR2_1416 (.Y(N4008),.A(N3951),.B(N3832));
NOR2X1 NOR2_1417 (.Y(N4009),.A(N3902),.B(N3955));
NOR2X1 NOR2_1418 (.Y(N4010),.A(N3955),.B(N3837));
NOR2X1 NOR2_1419 (.Y(N4011),.A(N3905),.B(N3959));
NOR2X1 NOR2_1420 (.Y(N4012),.A(N3959),.B(N3842));
NOR2X1 NOR2_1421 (.Y(N4013),.A(N3908),.B(N3963));
NOR2X1 NOR2_1422 (.Y(N4014),.A(N3963),.B(N3847));
NOR2X1 NOR2_1423 (.Y(N4015),.A(N3911),.B(N3967));
NOR2X1 NOR2_1424 (.Y(N4016),.A(N3967),.B(N3852));
NOR2X1 NOR2_1425 (.Y(N4017),.A(N3914),.B(N3971));
NOR2X1 NOR2_1426 (.Y(N4018),.A(N3971),.B(N3857));
NOR2X1 NOR2_1427 (.Y(N4019),.A(N3975),.B(N3976));
NOR2X1 NOR2_1428 (.Y(N4022),.A(N3977),.B(N954));
NOR2X1 NOR2_1429 (.Y(N4026),.A(N3923),.B(N3980));
NOR2X1 NOR2_1430 (.Y(N4027),.A(N3980),.B(N1002));
NOR2X1 NOR2_1431 (.Y(N4028),.A(N3800),.B(N3980));
NOR2X1 NOR2_1432 (.Y(N4031),.A(N3984),.B(N3985));
NOR2X1 NOR2_1433 (.Y(N4034),.A(N3989),.B(N3986));
NOR2X1 NOR2_1434 (.Y(N4038),.A(N3935),.B(N3992));
NOR2X1 NOR2_1435 (.Y(N4039),.A(N3992),.B(N3932));
NOR2X1 NOR2_1436 (.Y(N4040),.A(N3996),.B(N3997));
NOR2X1 NOR2_1437 (.Y(N4043),.A(N3998),.B(N1197));
NOR2X1 NOR2_1438 (.Y(N4047),.A(N3944),.B(N4001));
NOR2X1 NOR2_1439 (.Y(N4048),.A(N4001),.B(N1245));
NOR2X1 NOR2_1440 (.Y(N4049),.A(N3821),.B(N4001));
NOR2X1 NOR2_1441 (.Y(N4052),.A(N4005),.B(N4006));
NOR2X1 NOR2_1442 (.Y(N4055),.A(N4007),.B(N4008));
NOR2X1 NOR2_1443 (.Y(N4058),.A(N4009),.B(N4010));
NOR2X1 NOR2_1444 (.Y(N4061),.A(N4011),.B(N4012));
NOR2X1 NOR2_1445 (.Y(N4064),.A(N4013),.B(N4014));
NOR2X1 NOR2_1446 (.Y(N4067),.A(N4015),.B(N4016));
NOR2X1 NOR2_1447 (.Y(N4070),.A(N4017),.B(N4018));
NOR2X1 NOR2_1448 (.Y(N4073),.A(N4019),.B(N906));
NOR2X1 NOR2_1449 (.Y(N4077),.A(N3977),.B(N4022));
NOR2X1 NOR2_1450 (.Y(N4078),.A(N4022),.B(N954));
NOR2X1 NOR2_1451 (.Y(N4079),.A(N3868),.B(N4022));
NOR2X1 NOR2_1452 (.Y(N4082),.A(N4026),.B(N4027));
NOR2X1 NOR2_1453 (.Y(N4085),.A(N4031),.B(N4028));
NOR2X1 NOR2_1454 (.Y(N4089),.A(N3989),.B(N4034));
NOR2X1 NOR2_1455 (.Y(N4090),.A(N4034),.B(N3986));
NOR2X1 NOR2_1456 (.Y(N4091),.A(N4038),.B(N4039));
NOR2X1 NOR2_1457 (.Y(N4094),.A(N4040),.B(N1149));
NOR2X1 NOR2_1458 (.Y(N4098),.A(N3998),.B(N4043));
NOR2X1 NOR2_1459 (.Y(N4099),.A(N4043),.B(N1197));
NOR2X1 NOR2_1460 (.Y(N4100),.A(N3889),.B(N4043));
NOR2X1 NOR2_1461 (.Y(N4103),.A(N4047),.B(N4048));
NOR2X1 NOR2_1462 (.Y(N4106),.A(N1293),.B(N4049));
NOR2X1 NOR2_1463 (.Y(N4110),.A(N4052),.B(N570));
NOR2X1 NOR2_1464 (.Y(N4114),.A(N4055),.B(N618));
NOR2X1 NOR2_1465 (.Y(N4118),.A(N4058),.B(N666));
NOR2X1 NOR2_1466 (.Y(N4122),.A(N4061),.B(N714));
NOR2X1 NOR2_1467 (.Y(N4126),.A(N4064),.B(N762));
NOR2X1 NOR2_1468 (.Y(N4130),.A(N4067),.B(N810));
NOR2X1 NOR2_1469 (.Y(N4134),.A(N4070),.B(N858));
NOR2X1 NOR2_1470 (.Y(N4138),.A(N4019),.B(N4073));
NOR2X1 NOR2_1471 (.Y(N4139),.A(N4073),.B(N906));
NOR2X1 NOR2_1472 (.Y(N4140),.A(N3917),.B(N4073));
NOR2X1 NOR2_1473 (.Y(N4143),.A(N4077),.B(N4078));
NOR2X1 NOR2_1474 (.Y(N4146),.A(N4082),.B(N4079));
NOR2X1 NOR2_1475 (.Y(N4150),.A(N4031),.B(N4085));
NOR2X1 NOR2_1476 (.Y(N4151),.A(N4085),.B(N4028));
NOR2X1 NOR2_1477 (.Y(N4152),.A(N4089),.B(N4090));
NOR2X1 NOR2_1478 (.Y(N4155),.A(N4091),.B(N1101));
NOR2X1 NOR2_1479 (.Y(N4159),.A(N4040),.B(N4094));
NOR2X1 NOR2_1480 (.Y(N4160),.A(N4094),.B(N1149));
NOR2X1 NOR2_1481 (.Y(N4161),.A(N3938),.B(N4094));
NOR2X1 NOR2_1482 (.Y(N4164),.A(N4098),.B(N4099));
NOR2X1 NOR2_1483 (.Y(N4167),.A(N4103),.B(N4100));
NOR2X1 NOR2_1484 (.Y(N4171),.A(N1293),.B(N4106));
NOR2X1 NOR2_1485 (.Y(N4172),.A(N4106),.B(N4049));
NOR2X1 NOR2_1486 (.Y(N4173),.A(N4052),.B(N4110));
NOR2X1 NOR2_1487 (.Y(N4174),.A(N4110),.B(N570));
NOR2X1 NOR2_1488 (.Y(N4175),.A(N3947),.B(N4110));
NOR2X1 NOR2_1489 (.Y(N4178),.A(N4055),.B(N4114));
NOR2X1 NOR2_1490 (.Y(N4179),.A(N4114),.B(N618));
NOR2X1 NOR2_1491 (.Y(N4180),.A(N3951),.B(N4114));
NOR2X1 NOR2_1492 (.Y(N4183),.A(N4058),.B(N4118));
NOR2X1 NOR2_1493 (.Y(N4184),.A(N4118),.B(N666));
NOR2X1 NOR2_1494 (.Y(N4185),.A(N3955),.B(N4118));
NOR2X1 NOR2_1495 (.Y(N4188),.A(N4061),.B(N4122));
NOR2X1 NOR2_1496 (.Y(N4189),.A(N4122),.B(N714));
NOR2X1 NOR2_1497 (.Y(N4190),.A(N3959),.B(N4122));
NOR2X1 NOR2_1498 (.Y(N4193),.A(N4064),.B(N4126));
NOR2X1 NOR2_1499 (.Y(N4194),.A(N4126),.B(N762));
NOR2X1 NOR2_1500 (.Y(N4195),.A(N3963),.B(N4126));
NOR2X1 NOR2_1501 (.Y(N4198),.A(N4067),.B(N4130));
NOR2X1 NOR2_1502 (.Y(N4199),.A(N4130),.B(N810));
NOR2X1 NOR2_1503 (.Y(N4200),.A(N3967),.B(N4130));
NOR2X1 NOR2_1504 (.Y(N4203),.A(N4070),.B(N4134));
NOR2X1 NOR2_1505 (.Y(N4204),.A(N4134),.B(N858));
NOR2X1 NOR2_1506 (.Y(N4205),.A(N3971),.B(N4134));
NOR2X1 NOR2_1507 (.Y(N4208),.A(N4138),.B(N4139));
NOR2X1 NOR2_1508 (.Y(N4211),.A(N4143),.B(N4140));
NOR2X1 NOR2_1509 (.Y(N4215),.A(N4082),.B(N4146));
NOR2X1 NOR2_1510 (.Y(N4216),.A(N4146),.B(N4079));
NOR2X1 NOR2_1511 (.Y(N4217),.A(N4150),.B(N4151));
NOR2X1 NOR2_1512 (.Y(N4220),.A(N4152),.B(N1053));
NOR2X1 NOR2_1513 (.Y(N4224),.A(N4091),.B(N4155));
NOR2X1 NOR2_1514 (.Y(N4225),.A(N4155),.B(N1101));
NOR2X1 NOR2_1515 (.Y(N4226),.A(N3992),.B(N4155));
NOR2X1 NOR2_1516 (.Y(N4229),.A(N4159),.B(N4160));
NOR2X1 NOR2_1517 (.Y(N4232),.A(N4164),.B(N4161));
NOR2X1 NOR2_1518 (.Y(N4236),.A(N4103),.B(N4167));
NOR2X1 NOR2_1519 (.Y(N4237),.A(N4167),.B(N4100));
NOR2X1 NOR2_1520 (.Y(N4238),.A(N4171),.B(N4172));
NOR2X1 NOR2_1521 (.Y(N4241),.A(N4173),.B(N4174));
NOR2X1 NOR2_1522 (.Y(N4242),.A(N4178),.B(N4179));
NOR2X1 NOR2_1523 (.Y(N4245),.A(N4183),.B(N4184));
NOR2X1 NOR2_1524 (.Y(N4248),.A(N4188),.B(N4189));
NOR2X1 NOR2_1525 (.Y(N4251),.A(N4193),.B(N4194));
NOR2X1 NOR2_1526 (.Y(N4254),.A(N4198),.B(N4199));
NOR2X1 NOR2_1527 (.Y(N4257),.A(N4203),.B(N4204));
NOR2X1 NOR2_1528 (.Y(N4260),.A(N4208),.B(N4205));
NOR2X1 NOR2_1529 (.Y(N4264),.A(N4143),.B(N4211));
NOR2X1 NOR2_1530 (.Y(N4265),.A(N4211),.B(N4140));
NOR2X1 NOR2_1531 (.Y(N4266),.A(N4215),.B(N4216));
NOR2X1 NOR2_1532 (.Y(N4269),.A(N4217),.B(N1005));
NOR2X1 NOR2_1533 (.Y(N4273),.A(N4152),.B(N4220));
NOR2X1 NOR2_1534 (.Y(N4274),.A(N4220),.B(N1053));
NOR2X1 NOR2_1535 (.Y(N4275),.A(N4034),.B(N4220));
NOR2X1 NOR2_1536 (.Y(N4278),.A(N4224),.B(N4225));
NOR2X1 NOR2_1537 (.Y(N4281),.A(N4229),.B(N4226));
NOR2X1 NOR2_1538 (.Y(N4285),.A(N4164),.B(N4232));
NOR2X1 NOR2_1539 (.Y(N4286),.A(N4232),.B(N4161));
NOR2X1 NOR2_1540 (.Y(N4287),.A(N4236),.B(N4237));
NOR2X1 NOR2_1541 (.Y(N4290),.A(N4238),.B(N1248));
NOR2X1 NOR2_1542 (.Y(N4294),.A(N4242),.B(N4175));
NOR2X1 NOR2_1543 (.Y(N4298),.A(N4245),.B(N4180));
NOR2X1 NOR2_1544 (.Y(N4302),.A(N4248),.B(N4185));
NOR2X1 NOR2_1545 (.Y(N4306),.A(N4251),.B(N4190));
NOR2X1 NOR2_1546 (.Y(N4310),.A(N4254),.B(N4195));
NOR2X1 NOR2_1547 (.Y(N4314),.A(N4257),.B(N4200));
NOR2X1 NOR2_1548 (.Y(N4318),.A(N4208),.B(N4260));
NOR2X1 NOR2_1549 (.Y(N4319),.A(N4260),.B(N4205));
NOR2X1 NOR2_1550 (.Y(N4320),.A(N4264),.B(N4265));
NOR2X1 NOR2_1551 (.Y(N4323),.A(N4266),.B(N957));
NOR2X1 NOR2_1552 (.Y(N4327),.A(N4217),.B(N4269));
NOR2X1 NOR2_1553 (.Y(N4328),.A(N4269),.B(N1005));
NOR2X1 NOR2_1554 (.Y(N4329),.A(N4085),.B(N4269));
NOR2X1 NOR2_1555 (.Y(N4332),.A(N4273),.B(N4274));
NOR2X1 NOR2_1556 (.Y(N4335),.A(N4278),.B(N4275));
NOR2X1 NOR2_1557 (.Y(N4339),.A(N4229),.B(N4281));
NOR2X1 NOR2_1558 (.Y(N4340),.A(N4281),.B(N4226));
NOR2X1 NOR2_1559 (.Y(N4341),.A(N4285),.B(N4286));
NOR2X1 NOR2_1560 (.Y(N4344),.A(N4287),.B(N1200));
NOR2X1 NOR2_1561 (.Y(N4348),.A(N4238),.B(N4290));
NOR2X1 NOR2_1562 (.Y(N4349),.A(N4290),.B(N1248));
NOR2X1 NOR2_1563 (.Y(N4350),.A(N4106),.B(N4290));
NOR2X1 NOR2_1564 (.Y(N4353),.A(N4242),.B(N4294));
NOR2X1 NOR2_1565 (.Y(N4354),.A(N4294),.B(N4175));
NOR2X1 NOR2_1566 (.Y(N4355),.A(N4245),.B(N4298));
NOR2X1 NOR2_1567 (.Y(N4356),.A(N4298),.B(N4180));
NOR2X1 NOR2_1568 (.Y(N4357),.A(N4248),.B(N4302));
NOR2X1 NOR2_1569 (.Y(N4358),.A(N4302),.B(N4185));
NOR2X1 NOR2_1570 (.Y(N4359),.A(N4251),.B(N4306));
NOR2X1 NOR2_1571 (.Y(N4360),.A(N4306),.B(N4190));
NOR2X1 NOR2_1572 (.Y(N4361),.A(N4254),.B(N4310));
NOR2X1 NOR2_1573 (.Y(N4362),.A(N4310),.B(N4195));
NOR2X1 NOR2_1574 (.Y(N4363),.A(N4257),.B(N4314));
NOR2X1 NOR2_1575 (.Y(N4364),.A(N4314),.B(N4200));
NOR2X1 NOR2_1576 (.Y(N4365),.A(N4318),.B(N4319));
NOR2X1 NOR2_1577 (.Y(N4368),.A(N4320),.B(N909));
NOR2X1 NOR2_1578 (.Y(N4372),.A(N4266),.B(N4323));
NOR2X1 NOR2_1579 (.Y(N4373),.A(N4323),.B(N957));
NOR2X1 NOR2_1580 (.Y(N4374),.A(N4146),.B(N4323));
NOR2X1 NOR2_1581 (.Y(N4377),.A(N4327),.B(N4328));
NOR2X1 NOR2_1582 (.Y(N4380),.A(N4332),.B(N4329));
NOR2X1 NOR2_1583 (.Y(N4384),.A(N4278),.B(N4335));
NOR2X1 NOR2_1584 (.Y(N4385),.A(N4335),.B(N4275));
NOR2X1 NOR2_1585 (.Y(N4386),.A(N4339),.B(N4340));
NOR2X1 NOR2_1586 (.Y(N4389),.A(N4341),.B(N1152));
NOR2X1 NOR2_1587 (.Y(N4393),.A(N4287),.B(N4344));
NOR2X1 NOR2_1588 (.Y(N4394),.A(N4344),.B(N1200));
NOR2X1 NOR2_1589 (.Y(N4395),.A(N4167),.B(N4344));
NOR2X1 NOR2_1590 (.Y(N4398),.A(N4348),.B(N4349));
NOR2X1 NOR2_1591 (.Y(N4401),.A(N1296),.B(N4350));
NOR2X1 NOR2_1592 (.Y(N4405),.A(N4353),.B(N4354));
NOR2X1 NOR2_1593 (.Y(N4408),.A(N4355),.B(N4356));
NOR2X1 NOR2_1594 (.Y(N4411),.A(N4357),.B(N4358));
NOR2X1 NOR2_1595 (.Y(N4414),.A(N4359),.B(N4360));
NOR2X1 NOR2_1596 (.Y(N4417),.A(N4361),.B(N4362));
NOR2X1 NOR2_1597 (.Y(N4420),.A(N4363),.B(N4364));
NOR2X1 NOR2_1598 (.Y(N4423),.A(N4365),.B(N861));
NOR2X1 NOR2_1599 (.Y(N4427),.A(N4320),.B(N4368));
NOR2X1 NOR2_1600 (.Y(N4428),.A(N4368),.B(N909));
NOR2X1 NOR2_1601 (.Y(N4429),.A(N4211),.B(N4368));
NOR2X1 NOR2_1602 (.Y(N4432),.A(N4372),.B(N4373));
NOR2X1 NOR2_1603 (.Y(N4435),.A(N4377),.B(N4374));
NOR2X1 NOR2_1604 (.Y(N4439),.A(N4332),.B(N4380));
NOR2X1 NOR2_1605 (.Y(N4440),.A(N4380),.B(N4329));
NOR2X1 NOR2_1606 (.Y(N4441),.A(N4384),.B(N4385));
NOR2X1 NOR2_1607 (.Y(N4444),.A(N4386),.B(N1104));
NOR2X1 NOR2_1608 (.Y(N4448),.A(N4341),.B(N4389));
NOR2X1 NOR2_1609 (.Y(N4449),.A(N4389),.B(N1152));
NOR2X1 NOR2_1610 (.Y(N4450),.A(N4232),.B(N4389));
NOR2X1 NOR2_1611 (.Y(N4453),.A(N4393),.B(N4394));
NOR2X1 NOR2_1612 (.Y(N4456),.A(N4398),.B(N4395));
NOR2X1 NOR2_1613 (.Y(N4460),.A(N1296),.B(N4401));
NOR2X1 NOR2_1614 (.Y(N4461),.A(N4401),.B(N4350));
NOR2X1 NOR2_1615 (.Y(N4462),.A(N4405),.B(N573));
NOR2X1 NOR2_1616 (.Y(N4466),.A(N4408),.B(N621));
NOR2X1 NOR2_1617 (.Y(N4470),.A(N4411),.B(N669));
NOR2X1 NOR2_1618 (.Y(N4474),.A(N4414),.B(N717));
NOR2X1 NOR2_1619 (.Y(N4478),.A(N4417),.B(N765));
NOR2X1 NOR2_1620 (.Y(N4482),.A(N4420),.B(N813));
NOR2X1 NOR2_1621 (.Y(N4486),.A(N4365),.B(N4423));
NOR2X1 NOR2_1622 (.Y(N4487),.A(N4423),.B(N861));
NOR2X1 NOR2_1623 (.Y(N4488),.A(N4260),.B(N4423));
NOR2X1 NOR2_1624 (.Y(N4491),.A(N4427),.B(N4428));
NOR2X1 NOR2_1625 (.Y(N4494),.A(N4432),.B(N4429));
NOR2X1 NOR2_1626 (.Y(N4498),.A(N4377),.B(N4435));
NOR2X1 NOR2_1627 (.Y(N4499),.A(N4435),.B(N4374));
NOR2X1 NOR2_1628 (.Y(N4500),.A(N4439),.B(N4440));
NOR2X1 NOR2_1629 (.Y(N4503),.A(N4441),.B(N1056));
NOR2X1 NOR2_1630 (.Y(N4507),.A(N4386),.B(N4444));
NOR2X1 NOR2_1631 (.Y(N4508),.A(N4444),.B(N1104));
NOR2X1 NOR2_1632 (.Y(N4509),.A(N4281),.B(N4444));
NOR2X1 NOR2_1633 (.Y(N4512),.A(N4448),.B(N4449));
NOR2X1 NOR2_1634 (.Y(N4515),.A(N4453),.B(N4450));
NOR2X1 NOR2_1635 (.Y(N4519),.A(N4398),.B(N4456));
NOR2X1 NOR2_1636 (.Y(N4520),.A(N4456),.B(N4395));
NOR2X1 NOR2_1637 (.Y(N4521),.A(N4460),.B(N4461));
NOR2X1 NOR2_1638 (.Y(N4524),.A(N4405),.B(N4462));
NOR2X1 NOR2_1639 (.Y(N4525),.A(N4462),.B(N573));
NOR2X1 NOR2_1640 (.Y(N4526),.A(N4294),.B(N4462));
NOR2X1 NOR2_1641 (.Y(N4529),.A(N4408),.B(N4466));
NOR2X1 NOR2_1642 (.Y(N4530),.A(N4466),.B(N621));
NOR2X1 NOR2_1643 (.Y(N4531),.A(N4298),.B(N4466));
NOR2X1 NOR2_1644 (.Y(N4534),.A(N4411),.B(N4470));
NOR2X1 NOR2_1645 (.Y(N4535),.A(N4470),.B(N669));
NOR2X1 NOR2_1646 (.Y(N4536),.A(N4302),.B(N4470));
NOR2X1 NOR2_1647 (.Y(N4539),.A(N4414),.B(N4474));
NOR2X1 NOR2_1648 (.Y(N4540),.A(N4474),.B(N717));
NOR2X1 NOR2_1649 (.Y(N4541),.A(N4306),.B(N4474));
NOR2X1 NOR2_1650 (.Y(N4544),.A(N4417),.B(N4478));
NOR2X1 NOR2_1651 (.Y(N4545),.A(N4478),.B(N765));
NOR2X1 NOR2_1652 (.Y(N4546),.A(N4310),.B(N4478));
NOR2X1 NOR2_1653 (.Y(N4549),.A(N4420),.B(N4482));
NOR2X1 NOR2_1654 (.Y(N4550),.A(N4482),.B(N813));
NOR2X1 NOR2_1655 (.Y(N4551),.A(N4314),.B(N4482));
NOR2X1 NOR2_1656 (.Y(N4554),.A(N4486),.B(N4487));
NOR2X1 NOR2_1657 (.Y(N4557),.A(N4491),.B(N4488));
NOR2X1 NOR2_1658 (.Y(N4561),.A(N4432),.B(N4494));
NOR2X1 NOR2_1659 (.Y(N4562),.A(N4494),.B(N4429));
NOR2X1 NOR2_1660 (.Y(N4563),.A(N4498),.B(N4499));
NOR2X1 NOR2_1661 (.Y(N4566),.A(N4500),.B(N1008));
NOR2X1 NOR2_1662 (.Y(N4570),.A(N4441),.B(N4503));
NOR2X1 NOR2_1663 (.Y(N4571),.A(N4503),.B(N1056));
NOR2X1 NOR2_1664 (.Y(N4572),.A(N4335),.B(N4503));
NOR2X1 NOR2_1665 (.Y(N4575),.A(N4507),.B(N4508));
NOR2X1 NOR2_1666 (.Y(N4578),.A(N4512),.B(N4509));
NOR2X1 NOR2_1667 (.Y(N4582),.A(N4453),.B(N4515));
NOR2X1 NOR2_1668 (.Y(N4583),.A(N4515),.B(N4450));
NOR2X1 NOR2_1669 (.Y(N4584),.A(N4519),.B(N4520));
NOR2X1 NOR2_1670 (.Y(N4587),.A(N4521),.B(N1251));
NOR2X1 NOR2_1671 (.Y(N4591),.A(N4524),.B(N4525));
NOR2X1 NOR2_1672 (.Y(N4592),.A(N4529),.B(N4530));
NOR2X1 NOR2_1673 (.Y(N4595),.A(N4534),.B(N4535));
NOR2X1 NOR2_1674 (.Y(N4598),.A(N4539),.B(N4540));
NOR2X1 NOR2_1675 (.Y(N4601),.A(N4544),.B(N4545));
NOR2X1 NOR2_1676 (.Y(N4604),.A(N4549),.B(N4550));
NOR2X1 NOR2_1677 (.Y(N4607),.A(N4554),.B(N4551));
NOR2X1 NOR2_1678 (.Y(N4611),.A(N4491),.B(N4557));
NOR2X1 NOR2_1679 (.Y(N4612),.A(N4557),.B(N4488));
NOR2X1 NOR2_1680 (.Y(N4613),.A(N4561),.B(N4562));
NOR2X1 NOR2_1681 (.Y(N4616),.A(N4563),.B(N960));
NOR2X1 NOR2_1682 (.Y(N4620),.A(N4500),.B(N4566));
NOR2X1 NOR2_1683 (.Y(N4621),.A(N4566),.B(N1008));
NOR2X1 NOR2_1684 (.Y(N4622),.A(N4380),.B(N4566));
NOR2X1 NOR2_1685 (.Y(N4625),.A(N4570),.B(N4571));
NOR2X1 NOR2_1686 (.Y(N4628),.A(N4575),.B(N4572));
NOR2X1 NOR2_1687 (.Y(N4632),.A(N4512),.B(N4578));
NOR2X1 NOR2_1688 (.Y(N4633),.A(N4578),.B(N4509));
NOR2X1 NOR2_1689 (.Y(N4634),.A(N4582),.B(N4583));
NOR2X1 NOR2_1690 (.Y(N4637),.A(N4584),.B(N1203));
NOR2X1 NOR2_1691 (.Y(N4641),.A(N4521),.B(N4587));
NOR2X1 NOR2_1692 (.Y(N4642),.A(N4587),.B(N1251));
NOR2X1 NOR2_1693 (.Y(N4643),.A(N4401),.B(N4587));
NOR2X1 NOR2_1694 (.Y(N4646),.A(N4592),.B(N4526));
NOR2X1 NOR2_1695 (.Y(N4650),.A(N4595),.B(N4531));
NOR2X1 NOR2_1696 (.Y(N4654),.A(N4598),.B(N4536));
NOR2X1 NOR2_1697 (.Y(N4658),.A(N4601),.B(N4541));
NOR2X1 NOR2_1698 (.Y(N4662),.A(N4604),.B(N4546));
NOR2X1 NOR2_1699 (.Y(N4666),.A(N4554),.B(N4607));
NOR2X1 NOR2_1700 (.Y(N4667),.A(N4607),.B(N4551));
NOR2X1 NOR2_1701 (.Y(N4668),.A(N4611),.B(N4612));
NOR2X1 NOR2_1702 (.Y(N4671),.A(N4613),.B(N912));
NOR2X1 NOR2_1703 (.Y(N4675),.A(N4563),.B(N4616));
NOR2X1 NOR2_1704 (.Y(N4676),.A(N4616),.B(N960));
NOR2X1 NOR2_1705 (.Y(N4677),.A(N4435),.B(N4616));
NOR2X1 NOR2_1706 (.Y(N4680),.A(N4620),.B(N4621));
NOR2X1 NOR2_1707 (.Y(N4683),.A(N4625),.B(N4622));
NOR2X1 NOR2_1708 (.Y(N4687),.A(N4575),.B(N4628));
NOR2X1 NOR2_1709 (.Y(N4688),.A(N4628),.B(N4572));
NOR2X1 NOR2_1710 (.Y(N4689),.A(N4632),.B(N4633));
NOR2X1 NOR2_1711 (.Y(N4692),.A(N4634),.B(N1155));
NOR2X1 NOR2_1712 (.Y(N4696),.A(N4584),.B(N4637));
NOR2X1 NOR2_1713 (.Y(N4697),.A(N4637),.B(N1203));
NOR2X1 NOR2_1714 (.Y(N4698),.A(N4456),.B(N4637));
NOR2X1 NOR2_1715 (.Y(N4701),.A(N4641),.B(N4642));
NOR2X1 NOR2_1716 (.Y(N4704),.A(N1299),.B(N4643));
NOR2X1 NOR2_1717 (.Y(N4708),.A(N4592),.B(N4646));
NOR2X1 NOR2_1718 (.Y(N4709),.A(N4646),.B(N4526));
NOR2X1 NOR2_1719 (.Y(N4710),.A(N4595),.B(N4650));
NOR2X1 NOR2_1720 (.Y(N4711),.A(N4650),.B(N4531));
NOR2X1 NOR2_1721 (.Y(N4712),.A(N4598),.B(N4654));
NOR2X1 NOR2_1722 (.Y(N4713),.A(N4654),.B(N4536));
NOR2X1 NOR2_1723 (.Y(N4714),.A(N4601),.B(N4658));
NOR2X1 NOR2_1724 (.Y(N4715),.A(N4658),.B(N4541));
NOR2X1 NOR2_1725 (.Y(N4716),.A(N4604),.B(N4662));
NOR2X1 NOR2_1726 (.Y(N4717),.A(N4662),.B(N4546));
NOR2X1 NOR2_1727 (.Y(N4718),.A(N4666),.B(N4667));
NOR2X1 NOR2_1728 (.Y(N4721),.A(N4668),.B(N864));
NOR2X1 NOR2_1729 (.Y(N4725),.A(N4613),.B(N4671));
NOR2X1 NOR2_1730 (.Y(N4726),.A(N4671),.B(N912));
NOR2X1 NOR2_1731 (.Y(N4727),.A(N4494),.B(N4671));
NOR2X1 NOR2_1732 (.Y(N4730),.A(N4675),.B(N4676));
NOR2X1 NOR2_1733 (.Y(N4733),.A(N4680),.B(N4677));
NOR2X1 NOR2_1734 (.Y(N4737),.A(N4625),.B(N4683));
NOR2X1 NOR2_1735 (.Y(N4738),.A(N4683),.B(N4622));
NOR2X1 NOR2_1736 (.Y(N4739),.A(N4687),.B(N4688));
NOR2X1 NOR2_1737 (.Y(N4742),.A(N4689),.B(N1107));
NOR2X1 NOR2_1738 (.Y(N4746),.A(N4634),.B(N4692));
NOR2X1 NOR2_1739 (.Y(N4747),.A(N4692),.B(N1155));
NOR2X1 NOR2_1740 (.Y(N4748),.A(N4515),.B(N4692));
NOR2X1 NOR2_1741 (.Y(N4751),.A(N4696),.B(N4697));
NOR2X1 NOR2_1742 (.Y(N4754),.A(N4701),.B(N4698));
NOR2X1 NOR2_1743 (.Y(N4758),.A(N1299),.B(N4704));
NOR2X1 NOR2_1744 (.Y(N4759),.A(N4704),.B(N4643));
NOR2X1 NOR2_1745 (.Y(N4760),.A(N4708),.B(N4709));
NOR2X1 NOR2_1746 (.Y(N4763),.A(N4710),.B(N4711));
NOR2X1 NOR2_1747 (.Y(N4766),.A(N4712),.B(N4713));
NOR2X1 NOR2_1748 (.Y(N4769),.A(N4714),.B(N4715));
NOR2X1 NOR2_1749 (.Y(N4772),.A(N4716),.B(N4717));
NOR2X1 NOR2_1750 (.Y(N4775),.A(N4718),.B(N816));
NOR2X1 NOR2_1751 (.Y(N4779),.A(N4668),.B(N4721));
NOR2X1 NOR2_1752 (.Y(N4780),.A(N4721),.B(N864));
NOR2X1 NOR2_1753 (.Y(N4781),.A(N4557),.B(N4721));
NOR2X1 NOR2_1754 (.Y(N4784),.A(N4725),.B(N4726));
NOR2X1 NOR2_1755 (.Y(N4787),.A(N4730),.B(N4727));
NOR2X1 NOR2_1756 (.Y(N4791),.A(N4680),.B(N4733));
NOR2X1 NOR2_1757 (.Y(N4792),.A(N4733),.B(N4677));
NOR2X1 NOR2_1758 (.Y(N4793),.A(N4737),.B(N4738));
NOR2X1 NOR2_1759 (.Y(N4796),.A(N4739),.B(N1059));
NOR2X1 NOR2_1760 (.Y(N4800),.A(N4689),.B(N4742));
NOR2X1 NOR2_1761 (.Y(N4801),.A(N4742),.B(N1107));
NOR2X1 NOR2_1762 (.Y(N4802),.A(N4578),.B(N4742));
NOR2X1 NOR2_1763 (.Y(N4805),.A(N4746),.B(N4747));
NOR2X1 NOR2_1764 (.Y(N4808),.A(N4751),.B(N4748));
NOR2X1 NOR2_1765 (.Y(N4812),.A(N4701),.B(N4754));
NOR2X1 NOR2_1766 (.Y(N4813),.A(N4754),.B(N4698));
NOR2X1 NOR2_1767 (.Y(N4814),.A(N4758),.B(N4759));
NOR2X1 NOR2_1768 (.Y(N4817),.A(N4760),.B(N576));
NOR2X1 NOR2_1769 (.Y(N4821),.A(N4763),.B(N624));
NOR2X1 NOR2_1770 (.Y(N4825),.A(N4766),.B(N672));
NOR2X1 NOR2_1771 (.Y(N4829),.A(N4769),.B(N720));
NOR2X1 NOR2_1772 (.Y(N4833),.A(N4772),.B(N768));
NOR2X1 NOR2_1773 (.Y(N4837),.A(N4718),.B(N4775));
NOR2X1 NOR2_1774 (.Y(N4838),.A(N4775),.B(N816));
NOR2X1 NOR2_1775 (.Y(N4839),.A(N4607),.B(N4775));
NOR2X1 NOR2_1776 (.Y(N4842),.A(N4779),.B(N4780));
NOR2X1 NOR2_1777 (.Y(N4845),.A(N4784),.B(N4781));
NOR2X1 NOR2_1778 (.Y(N4849),.A(N4730),.B(N4787));
NOR2X1 NOR2_1779 (.Y(N4850),.A(N4787),.B(N4727));
NOR2X1 NOR2_1780 (.Y(N4851),.A(N4791),.B(N4792));
NOR2X1 NOR2_1781 (.Y(N4854),.A(N4793),.B(N1011));
NOR2X1 NOR2_1782 (.Y(N4858),.A(N4739),.B(N4796));
NOR2X1 NOR2_1783 (.Y(N4859),.A(N4796),.B(N1059));
NOR2X1 NOR2_1784 (.Y(N4860),.A(N4628),.B(N4796));
NOR2X1 NOR2_1785 (.Y(N4863),.A(N4800),.B(N4801));
NOR2X1 NOR2_1786 (.Y(N4866),.A(N4805),.B(N4802));
NOR2X1 NOR2_1787 (.Y(N4870),.A(N4751),.B(N4808));
NOR2X1 NOR2_1788 (.Y(N4871),.A(N4808),.B(N4748));
NOR2X1 NOR2_1789 (.Y(N4872),.A(N4812),.B(N4813));
NOR2X1 NOR2_1790 (.Y(N4875),.A(N4814),.B(N1254));
NOR2X1 NOR2_1791 (.Y(N4879),.A(N4760),.B(N4817));
NOR2X1 NOR2_1792 (.Y(N4880),.A(N4817),.B(N576));
NOR2X1 NOR2_1793 (.Y(N4881),.A(N4646),.B(N4817));
NOR2X1 NOR2_1794 (.Y(N4884),.A(N4763),.B(N4821));
NOR2X1 NOR2_1795 (.Y(N4885),.A(N4821),.B(N624));
NOR2X1 NOR2_1796 (.Y(N4886),.A(N4650),.B(N4821));
NOR2X1 NOR2_1797 (.Y(N4889),.A(N4766),.B(N4825));
NOR2X1 NOR2_1798 (.Y(N4890),.A(N4825),.B(N672));
NOR2X1 NOR2_1799 (.Y(N4891),.A(N4654),.B(N4825));
NOR2X1 NOR2_1800 (.Y(N4894),.A(N4769),.B(N4829));
NOR2X1 NOR2_1801 (.Y(N4895),.A(N4829),.B(N720));
NOR2X1 NOR2_1802 (.Y(N4896),.A(N4658),.B(N4829));
NOR2X1 NOR2_1803 (.Y(N4899),.A(N4772),.B(N4833));
NOR2X1 NOR2_1804 (.Y(N4900),.A(N4833),.B(N768));
NOR2X1 NOR2_1805 (.Y(N4901),.A(N4662),.B(N4833));
NOR2X1 NOR2_1806 (.Y(N4904),.A(N4837),.B(N4838));
NOR2X1 NOR2_1807 (.Y(N4907),.A(N4842),.B(N4839));
NOR2X1 NOR2_1808 (.Y(N4911),.A(N4784),.B(N4845));
NOR2X1 NOR2_1809 (.Y(N4912),.A(N4845),.B(N4781));
NOR2X1 NOR2_1810 (.Y(N4913),.A(N4849),.B(N4850));
NOR2X1 NOR2_1811 (.Y(N4916),.A(N4851),.B(N963));
NOR2X1 NOR2_1812 (.Y(N4920),.A(N4793),.B(N4854));
NOR2X1 NOR2_1813 (.Y(N4921),.A(N4854),.B(N1011));
NOR2X1 NOR2_1814 (.Y(N4922),.A(N4683),.B(N4854));
NOR2X1 NOR2_1815 (.Y(N4925),.A(N4858),.B(N4859));
NOR2X1 NOR2_1816 (.Y(N4928),.A(N4863),.B(N4860));
NOR2X1 NOR2_1817 (.Y(N4932),.A(N4805),.B(N4866));
NOR2X1 NOR2_1818 (.Y(N4933),.A(N4866),.B(N4802));
NOR2X1 NOR2_1819 (.Y(N4934),.A(N4870),.B(N4871));
NOR2X1 NOR2_1820 (.Y(N4937),.A(N4872),.B(N1206));
NOR2X1 NOR2_1821 (.Y(N4941),.A(N4814),.B(N4875));
NOR2X1 NOR2_1822 (.Y(N4942),.A(N4875),.B(N1254));
NOR2X1 NOR2_1823 (.Y(N4943),.A(N4704),.B(N4875));
NOR2X1 NOR2_1824 (.Y(N4946),.A(N4879),.B(N4880));
NOR2X1 NOR2_1825 (.Y(N4947),.A(N4884),.B(N4885));
NOR2X1 NOR2_1826 (.Y(N4950),.A(N4889),.B(N4890));
NOR2X1 NOR2_1827 (.Y(N4953),.A(N4894),.B(N4895));
NOR2X1 NOR2_1828 (.Y(N4956),.A(N4899),.B(N4900));
NOR2X1 NOR2_1829 (.Y(N4959),.A(N4904),.B(N4901));
NOR2X1 NOR2_1830 (.Y(N4963),.A(N4842),.B(N4907));
NOR2X1 NOR2_1831 (.Y(N4964),.A(N4907),.B(N4839));
NOR2X1 NOR2_1832 (.Y(N4965),.A(N4911),.B(N4912));
NOR2X1 NOR2_1833 (.Y(N4968),.A(N4913),.B(N915));
NOR2X1 NOR2_1834 (.Y(N4972),.A(N4851),.B(N4916));
NOR2X1 NOR2_1835 (.Y(N4973),.A(N4916),.B(N963));
NOR2X1 NOR2_1836 (.Y(N4974),.A(N4733),.B(N4916));
NOR2X1 NOR2_1837 (.Y(N4977),.A(N4920),.B(N4921));
NOR2X1 NOR2_1838 (.Y(N4980),.A(N4925),.B(N4922));
NOR2X1 NOR2_1839 (.Y(N4984),.A(N4863),.B(N4928));
NOR2X1 NOR2_1840 (.Y(N4985),.A(N4928),.B(N4860));
NOR2X1 NOR2_1841 (.Y(N4986),.A(N4932),.B(N4933));
NOR2X1 NOR2_1842 (.Y(N4989),.A(N4934),.B(N1158));
NOR2X1 NOR2_1843 (.Y(N4993),.A(N4872),.B(N4937));
NOR2X1 NOR2_1844 (.Y(N4994),.A(N4937),.B(N1206));
NOR2X1 NOR2_1845 (.Y(N4995),.A(N4754),.B(N4937));
NOR2X1 NOR2_1846 (.Y(N4998),.A(N4941),.B(N4942));
NOR2X1 NOR2_1847 (.Y(N5001),.A(N1302),.B(N4943));
NOR2X1 NOR2_1848 (.Y(N5005),.A(N4947),.B(N4881));
NOR2X1 NOR2_1849 (.Y(N5009),.A(N4950),.B(N4886));
NOR2X1 NOR2_1850 (.Y(N5013),.A(N4953),.B(N4891));
NOR2X1 NOR2_1851 (.Y(N5017),.A(N4956),.B(N4896));
NOR2X1 NOR2_1852 (.Y(N5021),.A(N4904),.B(N4959));
NOR2X1 NOR2_1853 (.Y(N5022),.A(N4959),.B(N4901));
NOR2X1 NOR2_1854 (.Y(N5023),.A(N4963),.B(N4964));
NOR2X1 NOR2_1855 (.Y(N5026),.A(N4965),.B(N867));
NOR2X1 NOR2_1856 (.Y(N5030),.A(N4913),.B(N4968));
NOR2X1 NOR2_1857 (.Y(N5031),.A(N4968),.B(N915));
NOR2X1 NOR2_1858 (.Y(N5032),.A(N4787),.B(N4968));
NOR2X1 NOR2_1859 (.Y(N5035),.A(N4972),.B(N4973));
NOR2X1 NOR2_1860 (.Y(N5038),.A(N4977),.B(N4974));
NOR2X1 NOR2_1861 (.Y(N5042),.A(N4925),.B(N4980));
NOR2X1 NOR2_1862 (.Y(N5043),.A(N4980),.B(N4922));
NOR2X1 NOR2_1863 (.Y(N5044),.A(N4984),.B(N4985));
NOR2X1 NOR2_1864 (.Y(N5047),.A(N4986),.B(N1110));
NOR2X1 NOR2_1865 (.Y(N5051),.A(N4934),.B(N4989));
NOR2X1 NOR2_1866 (.Y(N5052),.A(N4989),.B(N1158));
NOR2X1 NOR2_1867 (.Y(N5053),.A(N4808),.B(N4989));
NOR2X1 NOR2_1868 (.Y(N5056),.A(N4993),.B(N4994));
NOR2X1 NOR2_1869 (.Y(N5059),.A(N4998),.B(N4995));
NOR2X1 NOR2_1870 (.Y(N5063),.A(N1302),.B(N5001));
NOR2X1 NOR2_1871 (.Y(N5064),.A(N5001),.B(N4943));
NOR2X1 NOR2_1872 (.Y(N5065),.A(N4947),.B(N5005));
NOR2X1 NOR2_1873 (.Y(N5066),.A(N5005),.B(N4881));
NOR2X1 NOR2_1874 (.Y(N5067),.A(N4950),.B(N5009));
NOR2X1 NOR2_1875 (.Y(N5068),.A(N5009),.B(N4886));
NOR2X1 NOR2_1876 (.Y(N5069),.A(N4953),.B(N5013));
NOR2X1 NOR2_1877 (.Y(N5070),.A(N5013),.B(N4891));
NOR2X1 NOR2_1878 (.Y(N5071),.A(N4956),.B(N5017));
NOR2X1 NOR2_1879 (.Y(N5072),.A(N5017),.B(N4896));
NOR2X1 NOR2_1880 (.Y(N5073),.A(N5021),.B(N5022));
NOR2X1 NOR2_1881 (.Y(N5076),.A(N5023),.B(N819));
NOR2X1 NOR2_1882 (.Y(N5080),.A(N4965),.B(N5026));
NOR2X1 NOR2_1883 (.Y(N5081),.A(N5026),.B(N867));
NOR2X1 NOR2_1884 (.Y(N5082),.A(N4845),.B(N5026));
NOR2X1 NOR2_1885 (.Y(N5085),.A(N5030),.B(N5031));
NOR2X1 NOR2_1886 (.Y(N5088),.A(N5035),.B(N5032));
NOR2X1 NOR2_1887 (.Y(N5092),.A(N4977),.B(N5038));
NOR2X1 NOR2_1888 (.Y(N5093),.A(N5038),.B(N4974));
NOR2X1 NOR2_1889 (.Y(N5094),.A(N5042),.B(N5043));
NOR2X1 NOR2_1890 (.Y(N5097),.A(N5044),.B(N1062));
NOR2X1 NOR2_1891 (.Y(N5101),.A(N4986),.B(N5047));
NOR2X1 NOR2_1892 (.Y(N5102),.A(N5047),.B(N1110));
NOR2X1 NOR2_1893 (.Y(N5103),.A(N4866),.B(N5047));
NOR2X1 NOR2_1894 (.Y(N5106),.A(N5051),.B(N5052));
NOR2X1 NOR2_1895 (.Y(N5109),.A(N5056),.B(N5053));
NOR2X1 NOR2_1896 (.Y(N5113),.A(N4998),.B(N5059));
NOR2X1 NOR2_1897 (.Y(N5114),.A(N5059),.B(N4995));
NOR2X1 NOR2_1898 (.Y(N5115),.A(N5063),.B(N5064));
NOR2X1 NOR2_1899 (.Y(N5118),.A(N5065),.B(N5066));
NOR2X1 NOR2_1900 (.Y(N5121),.A(N5067),.B(N5068));
NOR2X1 NOR2_1901 (.Y(N5124),.A(N5069),.B(N5070));
NOR2X1 NOR2_1902 (.Y(N5127),.A(N5071),.B(N5072));
NOR2X1 NOR2_1903 (.Y(N5130),.A(N5073),.B(N771));
NOR2X1 NOR2_1904 (.Y(N5134),.A(N5023),.B(N5076));
NOR2X1 NOR2_1905 (.Y(N5135),.A(N5076),.B(N819));
NOR2X1 NOR2_1906 (.Y(N5136),.A(N4907),.B(N5076));
NOR2X1 NOR2_1907 (.Y(N5139),.A(N5080),.B(N5081));
NOR2X1 NOR2_1908 (.Y(N5142),.A(N5085),.B(N5082));
NOR2X1 NOR2_1909 (.Y(N5146),.A(N5035),.B(N5088));
NOR2X1 NOR2_1910 (.Y(N5147),.A(N5088),.B(N5032));
NOR2X1 NOR2_1911 (.Y(N5148),.A(N5092),.B(N5093));
NOR2X1 NOR2_1912 (.Y(N5151),.A(N5094),.B(N1014));
NOR2X1 NOR2_1913 (.Y(N5155),.A(N5044),.B(N5097));
NOR2X1 NOR2_1914 (.Y(N5156),.A(N5097),.B(N1062));
NOR2X1 NOR2_1915 (.Y(N5157),.A(N4928),.B(N5097));
NOR2X1 NOR2_1916 (.Y(N5160),.A(N5101),.B(N5102));
NOR2X1 NOR2_1917 (.Y(N5163),.A(N5106),.B(N5103));
NOR2X1 NOR2_1918 (.Y(N5167),.A(N5056),.B(N5109));
NOR2X1 NOR2_1919 (.Y(N5168),.A(N5109),.B(N5053));
NOR2X1 NOR2_1920 (.Y(N5169),.A(N5113),.B(N5114));
NOR2X1 NOR2_1921 (.Y(N5172),.A(N5115),.B(N1257));
NOR2X1 NOR2_1922 (.Y(N5176),.A(N5118),.B(N579));
NOR2X1 NOR2_1923 (.Y(N5180),.A(N5121),.B(N627));
NOR2X1 NOR2_1924 (.Y(N5184),.A(N5124),.B(N675));
NOR2X1 NOR2_1925 (.Y(N5188),.A(N5127),.B(N723));
NOR2X1 NOR2_1926 (.Y(N5192),.A(N5073),.B(N5130));
NOR2X1 NOR2_1927 (.Y(N5193),.A(N5130),.B(N771));
NOR2X1 NOR2_1928 (.Y(N5194),.A(N4959),.B(N5130));
NOR2X1 NOR2_1929 (.Y(N5197),.A(N5134),.B(N5135));
NOR2X1 NOR2_1930 (.Y(N5200),.A(N5139),.B(N5136));
NOR2X1 NOR2_1931 (.Y(N5204),.A(N5085),.B(N5142));
NOR2X1 NOR2_1932 (.Y(N5205),.A(N5142),.B(N5082));
NOR2X1 NOR2_1933 (.Y(N5206),.A(N5146),.B(N5147));
NOR2X1 NOR2_1934 (.Y(N5209),.A(N5148),.B(N966));
NOR2X1 NOR2_1935 (.Y(N5213),.A(N5094),.B(N5151));
NOR2X1 NOR2_1936 (.Y(N5214),.A(N5151),.B(N1014));
NOR2X1 NOR2_1937 (.Y(N5215),.A(N4980),.B(N5151));
NOR2X1 NOR2_1938 (.Y(N5218),.A(N5155),.B(N5156));
NOR2X1 NOR2_1939 (.Y(N5221),.A(N5160),.B(N5157));
NOR2X1 NOR2_1940 (.Y(N5225),.A(N5106),.B(N5163));
NOR2X1 NOR2_1941 (.Y(N5226),.A(N5163),.B(N5103));
NOR2X1 NOR2_1942 (.Y(N5227),.A(N5167),.B(N5168));
NOR2X1 NOR2_1943 (.Y(N5230),.A(N5169),.B(N1209));
NOR2X1 NOR2_1944 (.Y(N5234),.A(N5115),.B(N5172));
NOR2X1 NOR2_1945 (.Y(N5235),.A(N5172),.B(N1257));
NOR2X1 NOR2_1946 (.Y(N5236),.A(N5001),.B(N5172));
NOR2X1 NOR2_1947 (.Y(N5239),.A(N5118),.B(N5176));
NOR2X1 NOR2_1948 (.Y(N5240),.A(N5176),.B(N579));
NOR2X1 NOR2_1949 (.Y(N5241),.A(N5005),.B(N5176));
NOR2X1 NOR2_1950 (.Y(N5244),.A(N5121),.B(N5180));
NOR2X1 NOR2_1951 (.Y(N5245),.A(N5180),.B(N627));
NOR2X1 NOR2_1952 (.Y(N5246),.A(N5009),.B(N5180));
NOR2X1 NOR2_1953 (.Y(N5249),.A(N5124),.B(N5184));
NOR2X1 NOR2_1954 (.Y(N5250),.A(N5184),.B(N675));
NOR2X1 NOR2_1955 (.Y(N5251),.A(N5013),.B(N5184));
NOR2X1 NOR2_1956 (.Y(N5254),.A(N5127),.B(N5188));
NOR2X1 NOR2_1957 (.Y(N5255),.A(N5188),.B(N723));
NOR2X1 NOR2_1958 (.Y(N5256),.A(N5017),.B(N5188));
NOR2X1 NOR2_1959 (.Y(N5259),.A(N5192),.B(N5193));
NOR2X1 NOR2_1960 (.Y(N5262),.A(N5197),.B(N5194));
NOR2X1 NOR2_1961 (.Y(N5266),.A(N5139),.B(N5200));
NOR2X1 NOR2_1962 (.Y(N5267),.A(N5200),.B(N5136));
NOR2X1 NOR2_1963 (.Y(N5268),.A(N5204),.B(N5205));
NOR2X1 NOR2_1964 (.Y(N5271),.A(N5206),.B(N918));
NOR2X1 NOR2_1965 (.Y(N5275),.A(N5148),.B(N5209));
NOR2X1 NOR2_1966 (.Y(N5276),.A(N5209),.B(N966));
NOR2X1 NOR2_1967 (.Y(N5277),.A(N5038),.B(N5209));
NOR2X1 NOR2_1968 (.Y(N5280),.A(N5213),.B(N5214));
NOR2X1 NOR2_1969 (.Y(N5283),.A(N5218),.B(N5215));
NOR2X1 NOR2_1970 (.Y(N5287),.A(N5160),.B(N5221));
NOR2X1 NOR2_1971 (.Y(N5288),.A(N5221),.B(N5157));
NOR2X1 NOR2_1972 (.Y(N5289),.A(N5225),.B(N5226));
NOR2X1 NOR2_1973 (.Y(N5292),.A(N5227),.B(N1161));
NOR2X1 NOR2_1974 (.Y(N5296),.A(N5169),.B(N5230));
NOR2X1 NOR2_1975 (.Y(N5297),.A(N5230),.B(N1209));
NOR2X1 NOR2_1976 (.Y(N5298),.A(N5059),.B(N5230));
NOR2X1 NOR2_1977 (.Y(N5301),.A(N5234),.B(N5235));
NOR2X1 NOR2_1978 (.Y(N5304),.A(N1305),.B(N5236));
NOR2X1 NOR2_1979 (.Y(N5308),.A(N5239),.B(N5240));
NOR2X1 NOR2_1980 (.Y(N5309),.A(N5244),.B(N5245));
NOR2X1 NOR2_1981 (.Y(N5312),.A(N5249),.B(N5250));
NOR2X1 NOR2_1982 (.Y(N5315),.A(N5254),.B(N5255));
NOR2X1 NOR2_1983 (.Y(N5318),.A(N5259),.B(N5256));
NOR2X1 NOR2_1984 (.Y(N5322),.A(N5197),.B(N5262));
NOR2X1 NOR2_1985 (.Y(N5323),.A(N5262),.B(N5194));
NOR2X1 NOR2_1986 (.Y(N5324),.A(N5266),.B(N5267));
NOR2X1 NOR2_1987 (.Y(N5327),.A(N5268),.B(N870));
NOR2X1 NOR2_1988 (.Y(N5331),.A(N5206),.B(N5271));
NOR2X1 NOR2_1989 (.Y(N5332),.A(N5271),.B(N918));
NOR2X1 NOR2_1990 (.Y(N5333),.A(N5088),.B(N5271));
NOR2X1 NOR2_1991 (.Y(N5336),.A(N5275),.B(N5276));
NOR2X1 NOR2_1992 (.Y(N5339),.A(N5280),.B(N5277));
NOR2X1 NOR2_1993 (.Y(N5343),.A(N5218),.B(N5283));
NOR2X1 NOR2_1994 (.Y(N5344),.A(N5283),.B(N5215));
NOR2X1 NOR2_1995 (.Y(N5345),.A(N5287),.B(N5288));
NOR2X1 NOR2_1996 (.Y(N5348),.A(N5289),.B(N1113));
NOR2X1 NOR2_1997 (.Y(N5352),.A(N5227),.B(N5292));
NOR2X1 NOR2_1998 (.Y(N5353),.A(N5292),.B(N1161));
NOR2X1 NOR2_1999 (.Y(N5354),.A(N5109),.B(N5292));
NOR2X1 NOR2_2000 (.Y(N5357),.A(N5296),.B(N5297));
NOR2X1 NOR2_2001 (.Y(N5360),.A(N5301),.B(N5298));
NOR2X1 NOR2_2002 (.Y(N5364),.A(N1305),.B(N5304));
NOR2X1 NOR2_2003 (.Y(N5365),.A(N5304),.B(N5236));
NOR2X1 NOR2_2004 (.Y(N5366),.A(N5309),.B(N5241));
NOR2X1 NOR2_2005 (.Y(N5370),.A(N5312),.B(N5246));
NOR2X1 NOR2_2006 (.Y(N5374),.A(N5315),.B(N5251));
NOR2X1 NOR2_2007 (.Y(N5378),.A(N5259),.B(N5318));
NOR2X1 NOR2_2008 (.Y(N5379),.A(N5318),.B(N5256));
NOR2X1 NOR2_2009 (.Y(N5380),.A(N5322),.B(N5323));
NOR2X1 NOR2_2010 (.Y(N5383),.A(N5324),.B(N822));
NOR2X1 NOR2_2011 (.Y(N5387),.A(N5268),.B(N5327));
NOR2X1 NOR2_2012 (.Y(N5388),.A(N5327),.B(N870));
NOR2X1 NOR2_2013 (.Y(N5389),.A(N5142),.B(N5327));
NOR2X1 NOR2_2014 (.Y(N5392),.A(N5331),.B(N5332));
NOR2X1 NOR2_2015 (.Y(N5395),.A(N5336),.B(N5333));
NOR2X1 NOR2_2016 (.Y(N5399),.A(N5280),.B(N5339));
NOR2X1 NOR2_2017 (.Y(N5400),.A(N5339),.B(N5277));
NOR2X1 NOR2_2018 (.Y(N5401),.A(N5343),.B(N5344));
NOR2X1 NOR2_2019 (.Y(N5404),.A(N5345),.B(N1065));
NOR2X1 NOR2_2020 (.Y(N5408),.A(N5289),.B(N5348));
NOR2X1 NOR2_2021 (.Y(N5409),.A(N5348),.B(N1113));
NOR2X1 NOR2_2022 (.Y(N5410),.A(N5163),.B(N5348));
NOR2X1 NOR2_2023 (.Y(N5413),.A(N5352),.B(N5353));
NOR2X1 NOR2_2024 (.Y(N5416),.A(N5357),.B(N5354));
NOR2X1 NOR2_2025 (.Y(N5420),.A(N5301),.B(N5360));
NOR2X1 NOR2_2026 (.Y(N5421),.A(N5360),.B(N5298));
NOR2X1 NOR2_2027 (.Y(N5422),.A(N5364),.B(N5365));
NOR2X1 NOR2_2028 (.Y(N5425),.A(N5309),.B(N5366));
NOR2X1 NOR2_2029 (.Y(N5426),.A(N5366),.B(N5241));
NOR2X1 NOR2_2030 (.Y(N5427),.A(N5312),.B(N5370));
NOR2X1 NOR2_2031 (.Y(N5428),.A(N5370),.B(N5246));
NOR2X1 NOR2_2032 (.Y(N5429),.A(N5315),.B(N5374));
NOR2X1 NOR2_2033 (.Y(N5430),.A(N5374),.B(N5251));
NOR2X1 NOR2_2034 (.Y(N5431),.A(N5378),.B(N5379));
NOR2X1 NOR2_2035 (.Y(N5434),.A(N5380),.B(N774));
NOR2X1 NOR2_2036 (.Y(N5438),.A(N5324),.B(N5383));
NOR2X1 NOR2_2037 (.Y(N5439),.A(N5383),.B(N822));
NOR2X1 NOR2_2038 (.Y(N5440),.A(N5200),.B(N5383));
NOR2X1 NOR2_2039 (.Y(N5443),.A(N5387),.B(N5388));
NOR2X1 NOR2_2040 (.Y(N5446),.A(N5392),.B(N5389));
NOR2X1 NOR2_2041 (.Y(N5450),.A(N5336),.B(N5395));
NOR2X1 NOR2_2042 (.Y(N5451),.A(N5395),.B(N5333));
NOR2X1 NOR2_2043 (.Y(N5452),.A(N5399),.B(N5400));
NOR2X1 NOR2_2044 (.Y(N5455),.A(N5401),.B(N1017));
NOR2X1 NOR2_2045 (.Y(N5459),.A(N5345),.B(N5404));
NOR2X1 NOR2_2046 (.Y(N5460),.A(N5404),.B(N1065));
NOR2X1 NOR2_2047 (.Y(N5461),.A(N5221),.B(N5404));
NOR2X1 NOR2_2048 (.Y(N5464),.A(N5408),.B(N5409));
NOR2X1 NOR2_2049 (.Y(N5467),.A(N5413),.B(N5410));
NOR2X1 NOR2_2050 (.Y(N5471),.A(N5357),.B(N5416));
NOR2X1 NOR2_2051 (.Y(N5472),.A(N5416),.B(N5354));
NOR2X1 NOR2_2052 (.Y(N5473),.A(N5420),.B(N5421));
NOR2X1 NOR2_2053 (.Y(N5476),.A(N5422),.B(N1260));
NOR2X1 NOR2_2054 (.Y(N5480),.A(N5425),.B(N5426));
NOR2X1 NOR2_2055 (.Y(N5483),.A(N5427),.B(N5428));
NOR2X1 NOR2_2056 (.Y(N5486),.A(N5429),.B(N5430));
NOR2X1 NOR2_2057 (.Y(N5489),.A(N5431),.B(N726));
NOR2X1 NOR2_2058 (.Y(N5493),.A(N5380),.B(N5434));
NOR2X1 NOR2_2059 (.Y(N5494),.A(N5434),.B(N774));
NOR2X1 NOR2_2060 (.Y(N5495),.A(N5262),.B(N5434));
NOR2X1 NOR2_2061 (.Y(N5498),.A(N5438),.B(N5439));
NOR2X1 NOR2_2062 (.Y(N5501),.A(N5443),.B(N5440));
NOR2X1 NOR2_2063 (.Y(N5505),.A(N5392),.B(N5446));
NOR2X1 NOR2_2064 (.Y(N5506),.A(N5446),.B(N5389));
NOR2X1 NOR2_2065 (.Y(N5507),.A(N5450),.B(N5451));
NOR2X1 NOR2_2066 (.Y(N5510),.A(N5452),.B(N969));
NOR2X1 NOR2_2067 (.Y(N5514),.A(N5401),.B(N5455));
NOR2X1 NOR2_2068 (.Y(N5515),.A(N5455),.B(N1017));
NOR2X1 NOR2_2069 (.Y(N5516),.A(N5283),.B(N5455));
NOR2X1 NOR2_2070 (.Y(N5519),.A(N5459),.B(N5460));
NOR2X1 NOR2_2071 (.Y(N5522),.A(N5464),.B(N5461));
NOR2X1 NOR2_2072 (.Y(N5526),.A(N5413),.B(N5467));
NOR2X1 NOR2_2073 (.Y(N5527),.A(N5467),.B(N5410));
NOR2X1 NOR2_2074 (.Y(N5528),.A(N5471),.B(N5472));
NOR2X1 NOR2_2075 (.Y(N5531),.A(N5473),.B(N1212));
NOR2X1 NOR2_2076 (.Y(N5535),.A(N5422),.B(N5476));
NOR2X1 NOR2_2077 (.Y(N5536),.A(N5476),.B(N1260));
NOR2X1 NOR2_2078 (.Y(N5537),.A(N5304),.B(N5476));
NOR2X1 NOR2_2079 (.Y(N5540),.A(N5480),.B(N582));
NOR2X1 NOR2_2080 (.Y(N5544),.A(N5483),.B(N630));
NOR2X1 NOR2_2081 (.Y(N5548),.A(N5486),.B(N678));
NOR2X1 NOR2_2082 (.Y(N5552),.A(N5431),.B(N5489));
NOR2X1 NOR2_2083 (.Y(N5553),.A(N5489),.B(N726));
NOR2X1 NOR2_2084 (.Y(N5554),.A(N5318),.B(N5489));
NOR2X1 NOR2_2085 (.Y(N5557),.A(N5493),.B(N5494));
NOR2X1 NOR2_2086 (.Y(N5560),.A(N5498),.B(N5495));
NOR2X1 NOR2_2087 (.Y(N5564),.A(N5443),.B(N5501));
NOR2X1 NOR2_2088 (.Y(N5565),.A(N5501),.B(N5440));
NOR2X1 NOR2_2089 (.Y(N5566),.A(N5505),.B(N5506));
NOR2X1 NOR2_2090 (.Y(N5569),.A(N5507),.B(N921));
NOR2X1 NOR2_2091 (.Y(N5573),.A(N5452),.B(N5510));
NOR2X1 NOR2_2092 (.Y(N5574),.A(N5510),.B(N969));
NOR2X1 NOR2_2093 (.Y(N5575),.A(N5339),.B(N5510));
NOR2X1 NOR2_2094 (.Y(N5578),.A(N5514),.B(N5515));
NOR2X1 NOR2_2095 (.Y(N5581),.A(N5519),.B(N5516));
NOR2X1 NOR2_2096 (.Y(N5585),.A(N5464),.B(N5522));
NOR2X1 NOR2_2097 (.Y(N5586),.A(N5522),.B(N5461));
NOR2X1 NOR2_2098 (.Y(N5587),.A(N5526),.B(N5527));
NOR2X1 NOR2_2099 (.Y(N5590),.A(N5528),.B(N1164));
NOR2X1 NOR2_2100 (.Y(N5594),.A(N5473),.B(N5531));
NOR2X1 NOR2_2101 (.Y(N5595),.A(N5531),.B(N1212));
NOR2X1 NOR2_2102 (.Y(N5596),.A(N5360),.B(N5531));
NOR2X1 NOR2_2103 (.Y(N5599),.A(N5535),.B(N5536));
NOR2X1 NOR2_2104 (.Y(N5602),.A(N1308),.B(N5537));
NOR2X1 NOR2_2105 (.Y(N5606),.A(N5480),.B(N5540));
NOR2X1 NOR2_2106 (.Y(N5607),.A(N5540),.B(N582));
NOR2X1 NOR2_2107 (.Y(N5608),.A(N5366),.B(N5540));
NOR2X1 NOR2_2108 (.Y(N5611),.A(N5483),.B(N5544));
NOR2X1 NOR2_2109 (.Y(N5612),.A(N5544),.B(N630));
NOR2X1 NOR2_2110 (.Y(N5613),.A(N5370),.B(N5544));
NOR2X1 NOR2_2111 (.Y(N5616),.A(N5486),.B(N5548));
NOR2X1 NOR2_2112 (.Y(N5617),.A(N5548),.B(N678));
NOR2X1 NOR2_2113 (.Y(N5618),.A(N5374),.B(N5548));
NOR2X1 NOR2_2114 (.Y(N5621),.A(N5552),.B(N5553));
NOR2X1 NOR2_2115 (.Y(N5624),.A(N5557),.B(N5554));
NOR2X1 NOR2_2116 (.Y(N5628),.A(N5498),.B(N5560));
NOR2X1 NOR2_2117 (.Y(N5629),.A(N5560),.B(N5495));
NOR2X1 NOR2_2118 (.Y(N5630),.A(N5564),.B(N5565));
NOR2X1 NOR2_2119 (.Y(N5633),.A(N5566),.B(N873));
NOR2X1 NOR2_2120 (.Y(N5637),.A(N5507),.B(N5569));
NOR2X1 NOR2_2121 (.Y(N5638),.A(N5569),.B(N921));
NOR2X1 NOR2_2122 (.Y(N5639),.A(N5395),.B(N5569));
NOR2X1 NOR2_2123 (.Y(N5642),.A(N5573),.B(N5574));
NOR2X1 NOR2_2124 (.Y(N5645),.A(N5578),.B(N5575));
NOR2X1 NOR2_2125 (.Y(N5649),.A(N5519),.B(N5581));
NOR2X1 NOR2_2126 (.Y(N5650),.A(N5581),.B(N5516));
NOR2X1 NOR2_2127 (.Y(N5651),.A(N5585),.B(N5586));
NOR2X1 NOR2_2128 (.Y(N5654),.A(N5587),.B(N1116));
NOR2X1 NOR2_2129 (.Y(N5658),.A(N5528),.B(N5590));
NOR2X1 NOR2_2130 (.Y(N5659),.A(N5590),.B(N1164));
NOR2X1 NOR2_2131 (.Y(N5660),.A(N5416),.B(N5590));
NOR2X1 NOR2_2132 (.Y(N5663),.A(N5594),.B(N5595));
NOR2X1 NOR2_2133 (.Y(N5666),.A(N5599),.B(N5596));
NOR2X1 NOR2_2134 (.Y(N5670),.A(N1308),.B(N5602));
NOR2X1 NOR2_2135 (.Y(N5671),.A(N5602),.B(N5537));
NOR2X1 NOR2_2136 (.Y(N5672),.A(N5606),.B(N5607));
NOR2X1 NOR2_2137 (.Y(N5673),.A(N5611),.B(N5612));
NOR2X1 NOR2_2138 (.Y(N5676),.A(N5616),.B(N5617));
NOR2X1 NOR2_2139 (.Y(N5679),.A(N5621),.B(N5618));
NOR2X1 NOR2_2140 (.Y(N5683),.A(N5557),.B(N5624));
NOR2X1 NOR2_2141 (.Y(N5684),.A(N5624),.B(N5554));
NOR2X1 NOR2_2142 (.Y(N5685),.A(N5628),.B(N5629));
NOR2X1 NOR2_2143 (.Y(N5688),.A(N5630),.B(N825));
NOR2X1 NOR2_2144 (.Y(N5692),.A(N5566),.B(N5633));
NOR2X1 NOR2_2145 (.Y(N5693),.A(N5633),.B(N873));
NOR2X1 NOR2_2146 (.Y(N5694),.A(N5446),.B(N5633));
NOR2X1 NOR2_2147 (.Y(N5697),.A(N5637),.B(N5638));
NOR2X1 NOR2_2148 (.Y(N5700),.A(N5642),.B(N5639));
NOR2X1 NOR2_2149 (.Y(N5704),.A(N5578),.B(N5645));
NOR2X1 NOR2_2150 (.Y(N5705),.A(N5645),.B(N5575));
NOR2X1 NOR2_2151 (.Y(N5706),.A(N5649),.B(N5650));
NOR2X1 NOR2_2152 (.Y(N5709),.A(N5651),.B(N1068));
NOR2X1 NOR2_2153 (.Y(N5713),.A(N5587),.B(N5654));
NOR2X1 NOR2_2154 (.Y(N5714),.A(N5654),.B(N1116));
NOR2X1 NOR2_2155 (.Y(N5715),.A(N5467),.B(N5654));
NOR2X1 NOR2_2156 (.Y(N5718),.A(N5658),.B(N5659));
NOR2X1 NOR2_2157 (.Y(N5721),.A(N5663),.B(N5660));
NOR2X1 NOR2_2158 (.Y(N5725),.A(N5599),.B(N5666));
NOR2X1 NOR2_2159 (.Y(N5726),.A(N5666),.B(N5596));
NOR2X1 NOR2_2160 (.Y(N5727),.A(N5670),.B(N5671));
NOR2X1 NOR2_2161 (.Y(N5730),.A(N5673),.B(N5608));
NOR2X1 NOR2_2162 (.Y(N5734),.A(N5676),.B(N5613));
NOR2X1 NOR2_2163 (.Y(N5738),.A(N5621),.B(N5679));
NOR2X1 NOR2_2164 (.Y(N5739),.A(N5679),.B(N5618));
NOR2X1 NOR2_2165 (.Y(N5740),.A(N5683),.B(N5684));
NOR2X1 NOR2_2166 (.Y(N5743),.A(N5685),.B(N777));
NOR2X1 NOR2_2167 (.Y(N5747),.A(N5630),.B(N5688));
NOR2X1 NOR2_2168 (.Y(N5748),.A(N5688),.B(N825));
NOR2X1 NOR2_2169 (.Y(N5749),.A(N5501),.B(N5688));
NOR2X1 NOR2_2170 (.Y(N5752),.A(N5692),.B(N5693));
NOR2X1 NOR2_2171 (.Y(N5755),.A(N5697),.B(N5694));
NOR2X1 NOR2_2172 (.Y(N5759),.A(N5642),.B(N5700));
NOR2X1 NOR2_2173 (.Y(N5760),.A(N5700),.B(N5639));
NOR2X1 NOR2_2174 (.Y(N5761),.A(N5704),.B(N5705));
NOR2X1 NOR2_2175 (.Y(N5764),.A(N5706),.B(N1020));
NOR2X1 NOR2_2176 (.Y(N5768),.A(N5651),.B(N5709));
NOR2X1 NOR2_2177 (.Y(N5769),.A(N5709),.B(N1068));
NOR2X1 NOR2_2178 (.Y(N5770),.A(N5522),.B(N5709));
NOR2X1 NOR2_2179 (.Y(N5773),.A(N5713),.B(N5714));
NOR2X1 NOR2_2180 (.Y(N5776),.A(N5718),.B(N5715));
NOR2X1 NOR2_2181 (.Y(N5780),.A(N5663),.B(N5721));
NOR2X1 NOR2_2182 (.Y(N5781),.A(N5721),.B(N5660));
NOR2X1 NOR2_2183 (.Y(N5782),.A(N5725),.B(N5726));
NOR2X1 NOR2_2184 (.Y(N5785),.A(N5673),.B(N5730));
NOR2X1 NOR2_2185 (.Y(N5786),.A(N5730),.B(N5608));
NOR2X1 NOR2_2186 (.Y(N5787),.A(N5676),.B(N5734));
NOR2X1 NOR2_2187 (.Y(N5788),.A(N5734),.B(N5613));
NOR2X1 NOR2_2188 (.Y(N5789),.A(N5738),.B(N5739));
NOR2X1 NOR2_2189 (.Y(N5792),.A(N5740),.B(N729));
NOR2X1 NOR2_2190 (.Y(N5796),.A(N5685),.B(N5743));
NOR2X1 NOR2_2191 (.Y(N5797),.A(N5743),.B(N777));
NOR2X1 NOR2_2192 (.Y(N5798),.A(N5560),.B(N5743));
NOR2X1 NOR2_2193 (.Y(N5801),.A(N5747),.B(N5748));
NOR2X1 NOR2_2194 (.Y(N5804),.A(N5752),.B(N5749));
NOR2X1 NOR2_2195 (.Y(N5808),.A(N5697),.B(N5755));
NOR2X1 NOR2_2196 (.Y(N5809),.A(N5755),.B(N5694));
NOR2X1 NOR2_2197 (.Y(N5810),.A(N5759),.B(N5760));
NOR2X1 NOR2_2198 (.Y(N5813),.A(N5761),.B(N972));
NOR2X1 NOR2_2199 (.Y(N5817),.A(N5706),.B(N5764));
NOR2X1 NOR2_2200 (.Y(N5818),.A(N5764),.B(N1020));
NOR2X1 NOR2_2201 (.Y(N5819),.A(N5581),.B(N5764));
NOR2X1 NOR2_2202 (.Y(N5822),.A(N5768),.B(N5769));
NOR2X1 NOR2_2203 (.Y(N5825),.A(N5773),.B(N5770));
NOR2X1 NOR2_2204 (.Y(N5829),.A(N5718),.B(N5776));
NOR2X1 NOR2_2205 (.Y(N5830),.A(N5776),.B(N5715));
NOR2X1 NOR2_2206 (.Y(N5831),.A(N5780),.B(N5781));
NOR2X1 NOR2_2207 (.Y(N5834),.A(N5785),.B(N5786));
NOR2X1 NOR2_2208 (.Y(N5837),.A(N5787),.B(N5788));
NOR2X1 NOR2_2209 (.Y(N5840),.A(N5789),.B(N681));
NOR2X1 NOR2_2210 (.Y(N5844),.A(N5740),.B(N5792));
NOR2X1 NOR2_2211 (.Y(N5845),.A(N5792),.B(N729));
NOR2X1 NOR2_2212 (.Y(N5846),.A(N5624),.B(N5792));
NOR2X1 NOR2_2213 (.Y(N5849),.A(N5796),.B(N5797));
NOR2X1 NOR2_2214 (.Y(N5852),.A(N5801),.B(N5798));
NOR2X1 NOR2_2215 (.Y(N5856),.A(N5752),.B(N5804));
NOR2X1 NOR2_2216 (.Y(N5857),.A(N5804),.B(N5749));
NOR2X1 NOR2_2217 (.Y(N5858),.A(N5808),.B(N5809));
NOR2X1 NOR2_2218 (.Y(N5861),.A(N5810),.B(N924));
NOR2X1 NOR2_2219 (.Y(N5865),.A(N5761),.B(N5813));
NOR2X1 NOR2_2220 (.Y(N5866),.A(N5813),.B(N972));
NOR2X1 NOR2_2221 (.Y(N5867),.A(N5645),.B(N5813));
NOR2X1 NOR2_2222 (.Y(N5870),.A(N5817),.B(N5818));
NOR2X1 NOR2_2223 (.Y(N5873),.A(N5822),.B(N5819));
NOR2X1 NOR2_2224 (.Y(N5877),.A(N5773),.B(N5825));
NOR2X1 NOR2_2225 (.Y(N5878),.A(N5825),.B(N5770));
NOR2X1 NOR2_2226 (.Y(N5879),.A(N5829),.B(N5830));
NOR2X1 NOR2_2227 (.Y(N5882),.A(N5834),.B(N585));
NOR2X1 NOR2_2228 (.Y(N5886),.A(N5837),.B(N633));
NOR2X1 NOR2_2229 (.Y(N5890),.A(N5789),.B(N5840));
NOR2X1 NOR2_2230 (.Y(N5891),.A(N5840),.B(N681));
NOR2X1 NOR2_2231 (.Y(N5892),.A(N5679),.B(N5840));
NOR2X1 NOR2_2232 (.Y(N5895),.A(N5844),.B(N5845));
NOR2X1 NOR2_2233 (.Y(N5898),.A(N5849),.B(N5846));
NOR2X1 NOR2_2234 (.Y(N5902),.A(N5801),.B(N5852));
NOR2X1 NOR2_2235 (.Y(N5903),.A(N5852),.B(N5798));
NOR2X1 NOR2_2236 (.Y(N5904),.A(N5856),.B(N5857));
NOR2X1 NOR2_2237 (.Y(N5907),.A(N5858),.B(N876));
NOR2X1 NOR2_2238 (.Y(N5911),.A(N5810),.B(N5861));
NOR2X1 NOR2_2239 (.Y(N5912),.A(N5861),.B(N924));
NOR2X1 NOR2_2240 (.Y(N5913),.A(N5700),.B(N5861));
NOR2X1 NOR2_2241 (.Y(N5916),.A(N5865),.B(N5866));
NOR2X1 NOR2_2242 (.Y(N5919),.A(N5870),.B(N5867));
NOR2X1 NOR2_2243 (.Y(N5923),.A(N5822),.B(N5873));
NOR2X1 NOR2_2244 (.Y(N5924),.A(N5873),.B(N5819));
NOR2X1 NOR2_2245 (.Y(N5925),.A(N5877),.B(N5878));
NOR2X1 NOR2_2246 (.Y(N5928),.A(N5834),.B(N5882));
NOR2X1 NOR2_2247 (.Y(N5929),.A(N5882),.B(N585));
NOR2X1 NOR2_2248 (.Y(N5930),.A(N5730),.B(N5882));
NOR2X1 NOR2_2249 (.Y(N5933),.A(N5837),.B(N5886));
NOR2X1 NOR2_2250 (.Y(N5934),.A(N5886),.B(N633));
NOR2X1 NOR2_2251 (.Y(N5935),.A(N5734),.B(N5886));
NOR2X1 NOR2_2252 (.Y(N5938),.A(N5890),.B(N5891));
NOR2X1 NOR2_2253 (.Y(N5941),.A(N5895),.B(N5892));
NOR2X1 NOR2_2254 (.Y(N5945),.A(N5849),.B(N5898));
NOR2X1 NOR2_2255 (.Y(N5946),.A(N5898),.B(N5846));
NOR2X1 NOR2_2256 (.Y(N5947),.A(N5902),.B(N5903));
NOR2X1 NOR2_2257 (.Y(N5950),.A(N5904),.B(N828));
NOR2X1 NOR2_2258 (.Y(N5954),.A(N5858),.B(N5907));
NOR2X1 NOR2_2259 (.Y(N5955),.A(N5907),.B(N876));
NOR2X1 NOR2_2260 (.Y(N5956),.A(N5755),.B(N5907));
NOR2X1 NOR2_2261 (.Y(N5959),.A(N5911),.B(N5912));
NOR2X1 NOR2_2262 (.Y(N5962),.A(N5916),.B(N5913));
NOR2X1 NOR2_2263 (.Y(N5966),.A(N5870),.B(N5919));
NOR2X1 NOR2_2264 (.Y(N5967),.A(N5919),.B(N5867));
NOR2X1 NOR2_2265 (.Y(N5968),.A(N5923),.B(N5924));
NOR2X1 NOR2_2266 (.Y(N5971),.A(N5928),.B(N5929));
NOR2X1 NOR2_2267 (.Y(N5972),.A(N5933),.B(N5934));
NOR2X1 NOR2_2268 (.Y(N5975),.A(N5938),.B(N5935));
NOR2X1 NOR2_2269 (.Y(N5979),.A(N5895),.B(N5941));
NOR2X1 NOR2_2270 (.Y(N5980),.A(N5941),.B(N5892));
NOR2X1 NOR2_2271 (.Y(N5981),.A(N5945),.B(N5946));
NOR2X1 NOR2_2272 (.Y(N5984),.A(N5947),.B(N780));
NOR2X1 NOR2_2273 (.Y(N5988),.A(N5904),.B(N5950));
NOR2X1 NOR2_2274 (.Y(N5989),.A(N5950),.B(N828));
NOR2X1 NOR2_2275 (.Y(N5990),.A(N5804),.B(N5950));
NOR2X1 NOR2_2276 (.Y(N5993),.A(N5954),.B(N5955));
NOR2X1 NOR2_2277 (.Y(N5996),.A(N5959),.B(N5956));
NOR2X1 NOR2_2278 (.Y(N6000),.A(N5916),.B(N5962));
NOR2X1 NOR2_2279 (.Y(N6001),.A(N5962),.B(N5913));
NOR2X1 NOR2_2280 (.Y(N6002),.A(N5966),.B(N5967));
NOR2X1 NOR2_2281 (.Y(N6005),.A(N5972),.B(N5930));
NOR2X1 NOR2_2282 (.Y(N6009),.A(N5938),.B(N5975));
NOR2X1 NOR2_2283 (.Y(N6010),.A(N5975),.B(N5935));
NOR2X1 NOR2_2284 (.Y(N6011),.A(N5979),.B(N5980));
NOR2X1 NOR2_2285 (.Y(N6014),.A(N5981),.B(N732));
NOR2X1 NOR2_2286 (.Y(N6018),.A(N5947),.B(N5984));
NOR2X1 NOR2_2287 (.Y(N6019),.A(N5984),.B(N780));
NOR2X1 NOR2_2288 (.Y(N6020),.A(N5852),.B(N5984));
NOR2X1 NOR2_2289 (.Y(N6023),.A(N5988),.B(N5989));
NOR2X1 NOR2_2290 (.Y(N6026),.A(N5993),.B(N5990));
NOR2X1 NOR2_2291 (.Y(N6030),.A(N5959),.B(N5996));
NOR2X1 NOR2_2292 (.Y(N6031),.A(N5996),.B(N5956));
NOR2X1 NOR2_2293 (.Y(N6032),.A(N6000),.B(N6001));
NOR2X1 NOR2_2294 (.Y(N6035),.A(N5972),.B(N6005));
NOR2X1 NOR2_2295 (.Y(N6036),.A(N6005),.B(N5930));
NOR2X1 NOR2_2296 (.Y(N6037),.A(N6009),.B(N6010));
NOR2X1 NOR2_2297 (.Y(N6040),.A(N6011),.B(N684));
NOR2X1 NOR2_2298 (.Y(N6044),.A(N5981),.B(N6014));
NOR2X1 NOR2_2299 (.Y(N6045),.A(N6014),.B(N732));
NOR2X1 NOR2_2300 (.Y(N6046),.A(N5898),.B(N6014));
NOR2X1 NOR2_2301 (.Y(N6049),.A(N6018),.B(N6019));
NOR2X1 NOR2_2302 (.Y(N6052),.A(N6023),.B(N6020));
NOR2X1 NOR2_2303 (.Y(N6056),.A(N5993),.B(N6026));
NOR2X1 NOR2_2304 (.Y(N6057),.A(N6026),.B(N5990));
NOR2X1 NOR2_2305 (.Y(N6058),.A(N6030),.B(N6031));
NOR2X1 NOR2_2306 (.Y(N6061),.A(N6035),.B(N6036));
NOR2X1 NOR2_2307 (.Y(N6064),.A(N6037),.B(N636));
NOR2X1 NOR2_2308 (.Y(N6068),.A(N6011),.B(N6040));
NOR2X1 NOR2_2309 (.Y(N6069),.A(N6040),.B(N684));
NOR2X1 NOR2_2310 (.Y(N6070),.A(N5941),.B(N6040));
NOR2X1 NOR2_2311 (.Y(N6073),.A(N6044),.B(N6045));
NOR2X1 NOR2_2312 (.Y(N6076),.A(N6049),.B(N6046));
NOR2X1 NOR2_2313 (.Y(N6080),.A(N6023),.B(N6052));
NOR2X1 NOR2_2314 (.Y(N6081),.A(N6052),.B(N6020));
NOR2X1 NOR2_2315 (.Y(N6082),.A(N6056),.B(N6057));
NOR2X1 NOR2_2316 (.Y(N6085),.A(N6061),.B(N588));
NOR2X1 NOR2_2317 (.Y(N6089),.A(N6037),.B(N6064));
NOR2X1 NOR2_2318 (.Y(N6090),.A(N6064),.B(N636));
NOR2X1 NOR2_2319 (.Y(N6091),.A(N5975),.B(N6064));
NOR2X1 NOR2_2320 (.Y(N6094),.A(N6068),.B(N6069));
NOR2X1 NOR2_2321 (.Y(N6097),.A(N6073),.B(N6070));
NOR2X1 NOR2_2322 (.Y(N6101),.A(N6049),.B(N6076));
NOR2X1 NOR2_2323 (.Y(N6102),.A(N6076),.B(N6046));
NOR2X1 NOR2_2324 (.Y(N6103),.A(N6080),.B(N6081));
NOR2X1 NOR2_2325 (.Y(N6106),.A(N6061),.B(N6085));
NOR2X1 NOR2_2326 (.Y(N6107),.A(N6085),.B(N588));
NOR2X1 NOR2_2327 (.Y(N6108),.A(N6005),.B(N6085));
NOR2X1 NOR2_2328 (.Y(N6111),.A(N6089),.B(N6090));
NOR2X1 NOR2_2329 (.Y(N6114),.A(N6094),.B(N6091));
NOR2X1 NOR2_2330 (.Y(N6118),.A(N6073),.B(N6097));
NOR2X1 NOR2_2331 (.Y(N6119),.A(N6097),.B(N6070));
NOR2X1 NOR2_2332 (.Y(N6120),.A(N6101),.B(N6102));
NOR2X1 NOR2_2333 (.Y(N6123),.A(N6106),.B(N6107));
NOR2X1 NOR2_2334 (.Y(N6124),.A(N6111),.B(N6108));
NOR2X1 NOR2_2335 (.Y(N6128),.A(N6094),.B(N6114));
NOR2X1 NOR2_2336 (.Y(N6129),.A(N6114),.B(N6091));
NOR2X1 NOR2_2337 (.Y(N6130),.A(N6118),.B(N6119));
NOR2X1 NOR2_2338 (.Y(N6133),.A(N6111),.B(N6124));
NOR2X1 NOR2_2339 (.Y(N6134),.A(N6124),.B(N6108));
NOR2X1 NOR2_2340 (.Y(N6135),.A(N6128),.B(N6129));
NOR2X1 NOR2_2341 (.Y(N6138),.A(N6133),.B(N6134));
INVX1 NOT1_2342 (.Y(N6141),.A(N6138));
NOR2X1 NOR2_2343 (.Y(N6145),.A(N6138),.B(N6141));
INVX1 NOT1_2344 (.Y(N6146),.A(N6141));
NOR2X1 NOR2_2345 (.Y(N6147),.A(N6124),.B(N6141));
NOR2X1 NOR2_2346 (.Y(N6150),.A(N6145),.B(N6146));
NOR2X1 NOR2_2347 (.Y(N6151),.A(N6135),.B(N6147));
NOR2X1 NOR2_2348 (.Y(N6155),.A(N6135),.B(N6151));
NOR2X1 NOR2_2349 (.Y(N6156),.A(N6151),.B(N6147));
NOR2X1 NOR2_2350 (.Y(N6157),.A(N6114),.B(N6151));
NOR2X1 NOR2_2351 (.Y(N6160),.A(N6155),.B(N6156));
NOR2X1 NOR2_2352 (.Y(N6161),.A(N6130),.B(N6157));
NOR2X1 NOR2_2353 (.Y(N6165),.A(N6130),.B(N6161));
NOR2X1 NOR2_2354 (.Y(N6166),.A(N6161),.B(N6157));
NOR2X1 NOR2_2355 (.Y(N6167),.A(N6097),.B(N6161));
NOR2X1 NOR2_2356 (.Y(N6170),.A(N6165),.B(N6166));
NOR2X1 NOR2_2357 (.Y(N6171),.A(N6120),.B(N6167));
NOR2X1 NOR2_2358 (.Y(N6175),.A(N6120),.B(N6171));
NOR2X1 NOR2_2359 (.Y(N6176),.A(N6171),.B(N6167));
NOR2X1 NOR2_2360 (.Y(N6177),.A(N6076),.B(N6171));
NOR2X1 NOR2_2361 (.Y(N6180),.A(N6175),.B(N6176));
NOR2X1 NOR2_2362 (.Y(N6181),.A(N6103),.B(N6177));
NOR2X1 NOR2_2363 (.Y(N6185),.A(N6103),.B(N6181));
NOR2X1 NOR2_2364 (.Y(N6186),.A(N6181),.B(N6177));
NOR2X1 NOR2_2365 (.Y(N6187),.A(N6052),.B(N6181));
NOR2X1 NOR2_2366 (.Y(N6190),.A(N6185),.B(N6186));
NOR2X1 NOR2_2367 (.Y(N6191),.A(N6082),.B(N6187));
NOR2X1 NOR2_2368 (.Y(N6195),.A(N6082),.B(N6191));
NOR2X1 NOR2_2369 (.Y(N6196),.A(N6191),.B(N6187));
NOR2X1 NOR2_2370 (.Y(N6197),.A(N6026),.B(N6191));
NOR2X1 NOR2_2371 (.Y(N6200),.A(N6195),.B(N6196));
NOR2X1 NOR2_2372 (.Y(N6201),.A(N6058),.B(N6197));
NOR2X1 NOR2_2373 (.Y(N6205),.A(N6058),.B(N6201));
NOR2X1 NOR2_2374 (.Y(N6206),.A(N6201),.B(N6197));
NOR2X1 NOR2_2375 (.Y(N6207),.A(N5996),.B(N6201));
NOR2X1 NOR2_2376 (.Y(N6210),.A(N6205),.B(N6206));
NOR2X1 NOR2_2377 (.Y(N6211),.A(N6032),.B(N6207));
NOR2X1 NOR2_2378 (.Y(N6215),.A(N6032),.B(N6211));
NOR2X1 NOR2_2379 (.Y(N6216),.A(N6211),.B(N6207));
NOR2X1 NOR2_2380 (.Y(N6217),.A(N5962),.B(N6211));
NOR2X1 NOR2_2381 (.Y(N6220),.A(N6215),.B(N6216));
NOR2X1 NOR2_2382 (.Y(N6221),.A(N6002),.B(N6217));
NOR2X1 NOR2_2383 (.Y(N6225),.A(N6002),.B(N6221));
NOR2X1 NOR2_2384 (.Y(N6226),.A(N6221),.B(N6217));
NOR2X1 NOR2_2385 (.Y(N6227),.A(N5919),.B(N6221));
NOR2X1 NOR2_2386 (.Y(N6230),.A(N6225),.B(N6226));
NOR2X1 NOR2_2387 (.Y(N6231),.A(N5968),.B(N6227));
NOR2X1 NOR2_2388 (.Y(N6235),.A(N5968),.B(N6231));
NOR2X1 NOR2_2389 (.Y(N6236),.A(N6231),.B(N6227));
NOR2X1 NOR2_2390 (.Y(N6237),.A(N5873),.B(N6231));
NOR2X1 NOR2_2391 (.Y(N6240),.A(N6235),.B(N6236));
NOR2X1 NOR2_2392 (.Y(N6241),.A(N5925),.B(N6237));
NOR2X1 NOR2_2393 (.Y(N6245),.A(N5925),.B(N6241));
NOR2X1 NOR2_2394 (.Y(N6246),.A(N6241),.B(N6237));
NOR2X1 NOR2_2395 (.Y(N6247),.A(N5825),.B(N6241));
NOR2X1 NOR2_2396 (.Y(N6250),.A(N6245),.B(N6246));
NOR2X1 NOR2_2397 (.Y(N6251),.A(N5879),.B(N6247));
NOR2X1 NOR2_2398 (.Y(N6255),.A(N5879),.B(N6251));
NOR2X1 NOR2_2399 (.Y(N6256),.A(N6251),.B(N6247));
NOR2X1 NOR2_2400 (.Y(N6257),.A(N5776),.B(N6251));
NOR2X1 NOR2_2401 (.Y(N6260),.A(N6255),.B(N6256));
NOR2X1 NOR2_2402 (.Y(N6261),.A(N5831),.B(N6257));
NOR2X1 NOR2_2403 (.Y(N6265),.A(N5831),.B(N6261));
NOR2X1 NOR2_2404 (.Y(N6266),.A(N6261),.B(N6257));
NOR2X1 NOR2_2405 (.Y(N6267),.A(N5721),.B(N6261));
NOR2X1 NOR2_2406 (.Y(N6270),.A(N6265),.B(N6266));
NOR2X1 NOR2_2407 (.Y(N6271),.A(N5782),.B(N6267));
NOR2X1 NOR2_2408 (.Y(N6275),.A(N5782),.B(N6271));
NOR2X1 NOR2_2409 (.Y(N6276),.A(N6271),.B(N6267));
NOR2X1 NOR2_2410 (.Y(N6277),.A(N5666),.B(N6271));
NOR2X1 NOR2_2411 (.Y(N6280),.A(N6275),.B(N6276));
NOR2X1 NOR2_2412 (.Y(N6281),.A(N5727),.B(N6277));
NOR2X1 NOR2_2413 (.Y(N6285),.A(N5727),.B(N6281));
NOR2X1 NOR2_2414 (.Y(N6286),.A(N6281),.B(N6277));
NOR2X1 NOR2_2415 (.Y(N6287),.A(N5602),.B(N6281));
NOR2X1 NOR2_2416 (.Y(N6288),.A(N6285),.B(N6286));
endmodule 