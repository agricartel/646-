module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,N425,N428,N429;
INVX1 NOT1_1 (.Y(N118),.A(N1));
INVX1 NOT1_2 (.Y(N119),.A(N4));
INVX1 NOT1_3 (.Y(N122),.A(N11));
INVX1 NOT1_4 (.Y(N123),.A(N17));
INVX1 NOT1_5 (.Y(N126),.A(N24));
INVX1 NOT1_6 (.Y(N127),.A(N30));
INVX1 NOT1_7 (.Y(N130),.A(N37));
INVX1 NOT1_8 (.Y(N131),.A(N43));
INVX1 NOT1_9 (.Y(N134),.A(N50));
INVX1 NOT1_10 (.Y(N135),.A(N56));
INVX1 NOT1_11 (.Y(N138),.A(N63));
INVX1 NOT1_12 (.Y(N139),.A(N69));
INVX1 NOT1_13 (.Y(N142),.A(N76));
INVX1 NOT1_14 (.Y(N143),.A(N82));
INVX1 NOT1_15 (.Y(N146),.A(N89));
INVX1 NOT1_16 (.Y(N147),.A(N95));
INVX1 NOT1_17 (.Y(N150),.A(N102));
INVX1 NOT1_18 (.Y(N151),.A(N108));
NAND2X1 NAND2_19 (.Y(N154),.A(N118),.B(N4));
NOR2X1 NOR2_20 (.Y(N157),.A(N8),.B(N119));
NOR2X1 NOR2_21 (.Y(N158),.A(N14),.B(N119));
NAND2X1 NAND2_22 (.Y(N159),.A(N122),.B(N17));
NAND2X1 NAND2_23 (.Y(N162),.A(N126),.B(N30));
NAND2X1 NAND2_24 (.Y(N165),.A(N130),.B(N43));
NAND2X1 NAND2_25 (.Y(N168),.A(N134),.B(N56));
NAND2X1 NAND2_26 (.Y(N171),.A(N138),.B(N69));
NAND2X1 NAND2_27 (.Y(N174),.A(N142),.B(N82));
NAND2X1 NAND2_28 (.Y(N177),.A(N146),.B(N95));
NAND2X1 NAND2_29 (.Y(N180),.A(N150),.B(N108));
NOR2X1 NOR2_30 (.Y(N183),.A(N21),.B(N123));
NOR2X1 NOR2_31 (.Y(N184),.A(N27),.B(N123));
NOR2X1 NOR2_32 (.Y(N185),.A(N34),.B(N127));
NOR2X1 NOR2_33 (.Y(N186),.A(N40),.B(N127));
NOR2X1 NOR2_34 (.Y(N187),.A(N47),.B(N131));
NOR2X1 NOR2_35 (.Y(N188),.A(N53),.B(N131));
NOR2X1 NOR2_36 (.Y(N189),.A(N60),.B(N135));
NOR2X1 NOR2_37 (.Y(N190),.A(N66),.B(N135));
NOR2X1 NOR2_38 (.Y(N191),.A(N73),.B(N139));
NOR2X1 NOR2_39 (.Y(N192),.A(N79),.B(N139));
NOR2X1 NOR2_40 (.Y(N193),.A(N86),.B(N143));
NOR2X1 NOR2_41 (.Y(N194),.A(N92),.B(N143));
NOR2X1 NOR2_42 (.Y(N195),.A(N99),.B(N147));
NOR2X1 NOR2_43 (.Y(N196),.A(N105),.B(N147));
NOR2X1 NOR2_44 (.Y(N197),.A(N112),.B(N151));
NOR2X1 NOR2_45 (.Y(N198),.A(N115),.B(N151));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N177),.B(N180));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N154),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(ttmp3),.A(N159),.B(ttmp2));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N162),.B(ttmp3));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N165),.B(ttmp4));
AND2X1 AND_tmp6 (.Y(ttmp6),.A(N168),.B(ttmp5));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N171),.B(ttmp6));
AND2X1 AND_tmp8 (.Y(N199),.A(N174),.B(ttmp7));
INVX1 NOT1_47 (.Y(N203),.A(N199));
INVX1 NOT1_48 (.Y(N213),.A(N199));
INVX1 NOT1_49 (.Y(N223),.A(N199));
XOR2X1 XOR2_50 (.Y(N224),.A(N203),.B(N154));
XOR2X1 XOR2_51 (.Y(N227),.A(N203),.B(N159));
XOR2X1 XOR2_52 (.Y(N230),.A(N203),.B(N162));
XOR2X1 XOR2_53 (.Y(N233),.A(N203),.B(N165));
XOR2X1 XOR2_54 (.Y(N236),.A(N203),.B(N168));
XOR2X1 XOR2_55 (.Y(N239),.A(N203),.B(N171));
NAND2X1 NAND2_56 (.Y(N242),.A(N1),.B(N213));
XOR2X1 XOR2_57 (.Y(N243),.A(N203),.B(N174));
NAND2X1 NAND2_58 (.Y(N246),.A(N213),.B(N11));
XOR2X1 XOR2_59 (.Y(N247),.A(N203),.B(N177));
NAND2X1 NAND2_60 (.Y(N250),.A(N213),.B(N24));
XOR2X1 XOR2_61 (.Y(N251),.A(N203),.B(N180));
NAND2X1 NAND2_62 (.Y(N254),.A(N213),.B(N37));
NAND2X1 NAND2_63 (.Y(N255),.A(N213),.B(N50));
NAND2X1 NAND2_64 (.Y(N256),.A(N213),.B(N63));
NAND2X1 NAND2_65 (.Y(N257),.A(N213),.B(N76));
NAND2X1 NAND2_66 (.Y(N258),.A(N213),.B(N89));
NAND2X1 NAND2_67 (.Y(N259),.A(N213),.B(N102));
NAND2X1 NAND2_68 (.Y(N260),.A(N224),.B(N157));
NAND2X1 NAND2_69 (.Y(N263),.A(N224),.B(N158));
NAND2X1 NAND2_70 (.Y(N264),.A(N227),.B(N183));
NAND2X1 NAND2_71 (.Y(N267),.A(N230),.B(N185));
NAND2X1 NAND2_72 (.Y(N270),.A(N233),.B(N187));
NAND2X1 NAND2_73 (.Y(N273),.A(N236),.B(N189));
AND2X1 NAND2_74 (.Y(N276),.A(N239),.B(N191));
NAND2X1 NAND2_75 (.Y(N279),.A(N243),.B(N193));
NAND2X1 NAND2_76 (.Y(N282),.A(N247),.B(N195));
NAND2X1 NAND2_77 (.Y(N285),.A(N251),.B(N197));
NAND2X1 NAND2_78 (.Y(N288),.A(N227),.B(N184));
NAND2X1 NAND2_79 (.Y(N289),.A(N230),.B(N186));
NAND2X1 NAND2_80 (.Y(N290),.A(N233),.B(N188));
NAND2X1 NAND2_81 (.Y(N291),.A(N236),.B(N190));
NAND2X1 NAND2_82 (.Y(N292),.A(N239),.B(N192));
NAND2X1 NAND2_83 (.Y(N293),.A(N243),.B(N194));
NAND2X1 NAND2_84 (.Y(N294),.A(N247),.B(N196));
NAND2X1 NAND2_85 (.Y(N295),.A(N251),.B(N198));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(N282),.B(N285));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N260),.B(ttmp9));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(N264),.B(ttmp10));
XOR2X1 AND_tmp12 (.Y(ttmp12),.A(N267),.B(ttmp11));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(N270),.B(ttmp12));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(N273),.B(ttmp13));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(N276),.B(ttmp14));
AND2X1 AND_tmp16 (.Y(N296),.A(N279),.B(ttmp15));
INVX1 NOT1_87 (.Y(N300),.A(N263));
INVX1 NOT1_88 (.Y(N301),.A(N288));
INVX1 NOT1_89 (.Y(N302),.A(N289));
INVX1 NOT1_90 (.Y(N303),.A(N290));
INVX1 NOT1_91 (.Y(N304),.A(N291));
INVX1 NOT1_92 (.Y(N305),.A(N292));
INVX1 NOT1_93 (.Y(N306),.A(N293));
INVX1 NOT1_94 (.Y(N307),.A(N294));
INVX1 NOT1_95 (.Y(N308),.A(N295));
INVX1 NOT1_96 (.Y(N309),.A(N296));
INVX1 NOT1_97 (.Y(N319),.A(N296));
INVX1 NOT1_98 (.Y(N329),.A(N296));
XOR2X1 XOR2_99 (.Y(N330),.A(N309),.B(N260));
XOR2X1 XOR2_100 (.Y(N331),.A(N309),.B(N264));
XOR2X1 XOR2_101 (.Y(N332),.A(N309),.B(N267));
XOR2X1 XOR2_102 (.Y(N333),.A(N309),.B(N270));
NAND2X1 NAND2_103 (.Y(N334),.A(N8),.B(N319));
XOR2X1 XOR2_104 (.Y(N335),.A(N309),.B(N273));
NAND2X1 NAND2_105 (.Y(N336),.A(N319),.B(N21));
XOR2X1 XOR2_106 (.Y(N337),.A(N309),.B(N276));
NAND2X1 NAND2_107 (.Y(N338),.A(N319),.B(N34));
XOR2X1 XOR2_108 (.Y(N339),.A(N309),.B(N279));
NAND2X1 NAND2_109 (.Y(N340),.A(N319),.B(N47));
XOR2X1 XOR2_110 (.Y(N341),.A(N309),.B(N282));
NAND2X1 NAND2_111 (.Y(N342),.A(N319),.B(N60));
XOR2X1 XOR2_112 (.Y(N343),.A(N309),.B(N285));
NAND2X1 NAND2_113 (.Y(N344),.A(N319),.B(N73));
NAND2X1 NAND2_114 (.Y(N345),.A(N319),.B(N86));
NAND2X1 NAND2_115 (.Y(N346),.A(N319),.B(N99));
NAND2X1 NAND2_116 (.Y(N347),.A(N319),.B(N112));
NAND2X1 NAND2_117 (.Y(N348),.A(N330),.B(N300));
NAND2X1 NAND2_118 (.Y(N349),.A(N331),.B(N301));
NAND2X1 NAND2_119 (.Y(N350),.A(N332),.B(N302));
NAND2X1 NAND2_120 (.Y(N351),.A(N333),.B(N303));
NAND2X1 NAND2_121 (.Y(N352),.A(N335),.B(N304));
NAND2X1 NAND2_122 (.Y(N353),.A(N337),.B(N305));
NAND2X1 NAND2_123 (.Y(N354),.A(N339),.B(N306));
NAND2X1 NAND2_124 (.Y(N355),.A(N341),.B(N307));
NAND2X1 NAND2_125 (.Y(N356),.A(N343),.B(N308));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N355),.B(N356));
AND2X1 AND_tmp18 (.Y(ttmp18),.A(N348),.B(ttmp17));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(N349),.B(ttmp18));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N350),.B(ttmp19));
AND2X1 AND_tmp21 (.Y(ttmp21),.A(N351),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N352),.B(ttmp21));
AND2X1 AND_tmp23 (.Y(ttmp23),.A(N353),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(N357),.A(N354),.B(ttmp23));
INVX1 NOT1_127 (.Y(N360),.A(N357));
INVX1 NOT1_128 (.Y(N370),.A(N357));
NAND2X1 NAND2_129 (.Y(N371),.A(N14),.B(N360));
NAND2X1 NAND2_130 (.Y(N372),.A(N360),.B(N27));
NAND2X1 NAND2_131 (.Y(N373),.A(N360),.B(N40));
NAND2X1 NAND2_132 (.Y(N374),.A(N360),.B(N53));
NAND2X1 NAND2_133 (.Y(N375),.A(N360),.B(N66));
NAND2X1 NAND2_134 (.Y(N376),.A(N360),.B(N79));
NAND2X1 NAND2_135 (.Y(N377),.A(N360),.B(N92));
NAND2X1 NAND2_136 (.Y(N378),.A(N360),.B(N105));
NAND2X1 NAND2_137 (.Y(N379),.A(N360),.B(N115));
AND2X1 AND_tmp25 (.Y(ttmp25),.A(N334),.B(N371));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N4),.B(ttmp25));
NAND2X1 NAND_tmp27 (.Y(N380),.A(N242),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(ttmp28),.A(N372),.B(N17));
AND2X1 AND_tmp29 (.Y(ttmp29),.A(N246),.B(ttmp28));
NAND2X1 NAND_tmp30 (.Y(N381),.A(N336),.B(ttmp29));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(N373),.B(N30));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(N250),.B(ttmp31));
NAND2X1 NAND_tmp33 (.Y(N386),.A(N338),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N374),.B(N43));
AND2X1 AND_tmp35 (.Y(ttmp35),.A(N254),.B(ttmp34));
NAND2X1 NAND_tmp36 (.Y(N393),.A(N340),.B(ttmp35));
AND2X1 AND_tmp37 (.Y(ttmp37),.A(N375),.B(N56));
XOR2X1 AND_tmp38 (.Y(ttmp38),.A(N255),.B(ttmp37));
NAND2X1 NAND_tmp39 (.Y(N399),.A(N342),.B(ttmp38));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N376),.B(N69));
AND2X1 AND_tmp41 (.Y(ttmp41),.A(N256),.B(ttmp40));
NAND2X1 NAND_tmp42 (.Y(N404),.A(N344),.B(ttmp41));
AND2X1 AND_tmp43 (.Y(ttmp43),.A(N377),.B(N82));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N257),.B(ttmp43));
NAND2X1 NAND_tmp45 (.Y(N407),.A(N345),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(N378),.B(N95));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(N258),.B(ttmp46));
NAND2X1 NAND_tmp48 (.Y(N411),.A(N346),.B(ttmp47));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(N379),.B(N108));
AND2X1 AND_tmp50 (.Y(ttmp50),.A(N259),.B(ttmp49));
NAND2X1 NAND_tmp51 (.Y(N414),.A(N347),.B(ttmp50));
INVX1 NOT1_147 (.Y(N415),.A(N380));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(N411),.B(N414));
AND2X1 AND_tmp53 (.Y(ttmp53),.A(N381),.B(ttmp52));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N386),.B(ttmp53));
AND2X1 AND_tmp55 (.Y(ttmp55),.A(N393),.B(ttmp54));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N399),.B(ttmp55));
AND2X1 AND_tmp57 (.Y(ttmp57),.A(N404),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(N416),.A(N407),.B(ttmp57));
INVX1 NOT1_149 (.Y(N417),.A(N393));
INVX1 NOT1_150 (.Y(N418),.A(N404));
INVX1 NOT1_151 (.Y(N419),.A(N407));
INVX1 NOT1_152 (.Y(N420),.A(N411));
NOR2X1 NOR2_153 (.Y(N421),.A(N415),.B(N416));
NAND2X1 NAND2_154 (.Y(N422),.A(N386),.B(N417));
AND2X1 AND_tmp59 (.Y(ttmp59),.A(N418),.B(N399));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N386),.B(ttmp59));
NAND2X1 NAND_tmp61 (.Y(N425),.A(N393),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N393),.B(N419));
NAND2X1 NAND_tmp63 (.Y(N428),.A(N399),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(ttmp64),.A(N407),.B(N420));
AND2X1 AND_tmp65 (.Y(ttmp65),.A(N386),.B(ttmp64));
NAND2X1 NAND_tmp66 (.Y(N429),.A(N393),.B(ttmp65));
AND2X1 AND_tmp67 (.Y(ttmp67),.A(N422),.B(N399));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N381),.B(ttmp67));
NAND2X1 NAND_tmp69 (.Y(N430),.A(N386),.B(ttmp68));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N425),.B(N428));
AND2X1 AND_tmp71 (.Y(ttmp71),.A(N381),.B(ttmp70));
NAND2X1 NAND_tmp72 (.Y(N431),.A(N386),.B(ttmp71));
AND2X1 AND_tmp73 (.Y(ttmp73),.A(N425),.B(N429));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N381),.B(ttmp73));
NAND2X1 NAND_tmp75 (.Y(N432),.A(N422),.B(ttmp74));
endmodule 