module c1355 (G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;
wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,G284,G287,G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,G329,G332,G335,G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,G421,G422,G423,G424,G425,G426,G429,G432,G435,G438,G441,G444,G447,G450,G453,G456,G459,G462,G465,G468,G471,G474,G477,G480,G483,G486,G489,G492,G495,G498,G501,G504,G507,G510,G513,G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,G546,G549,G552,G555,G558,G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,G642,G645,G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,G751,G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,G809,G812,G815,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,G986,G991,G996,G1001,G1006,G1011,G1016,G1021,G1026,G1031,G1036,G1039,G1042,G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,G1078,G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,G1117,G1120,G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,G1153,G1156,G1159,G1162,G1165,G1168,G1171,G1174,G1177,G1180,G1183,G1186,G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,G1222,G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,G1322,G1323;
AND2X1 AND2_0 (.Y(G242),.A(G33),.B(G41));
AND2X1 AND2_1 (.Y(G245),.A(G34),.B(G41));
AND2X1 AND2_2 (.Y(G248),.A(G35),.B(G41));
AND2X1 AND2_3 (.Y(G251),.A(G36),.B(G41));
AND2X1 AND2_4 (.Y(G254),.A(G37),.B(G41));
AND2X1 AND2_5 (.Y(G257),.A(G38),.B(G41));
AND2X1 AND2_6 (.Y(G260),.A(G39),.B(G41));
AND2X1 AND2_7 (.Y(G263),.A(G40),.B(G41));
NAND2X1 NAND2_0 (.Y(G266),.A(G1),.B(G2));
NAND2X1 NAND2_1 (.Y(G269),.A(G3),.B(G4));
NAND2X1 NAND2_2 (.Y(G272),.A(G5),.B(G6));
NAND2X1 NAND2_3 (.Y(G275),.A(G7),.B(G8));
NAND2X1 NAND2_4 (.Y(G278),.A(G9),.B(G10));
NAND2X1 NAND2_5 (.Y(G281),.A(G11),.B(G12));
NAND2X1 NAND2_6 (.Y(G284),.A(G13),.B(G14));
NAND2X1 NAND2_7 (.Y(G287),.A(G15),.B(G16));
NAND2X1 NAND2_8 (.Y(G290),.A(G17),.B(G18));
NAND2X1 NAND2_9 (.Y(G293),.A(G19),.B(G20));
NAND2X1 NAND2_10 (.Y(G296),.A(G21),.B(G22));
NAND2X1 NAND2_11 (.Y(G299),.A(G23),.B(G24));
NAND2X1 NAND2_12 (.Y(G302),.A(G25),.B(G26));
NAND2X1 NAND2_13 (.Y(G305),.A(G27),.B(G28));
NAND2X1 NAND2_14 (.Y(G308),.A(G29),.B(G30));
NAND2X1 NAND2_15 (.Y(G311),.A(G31),.B(G32));
NAND2X1 NAND2_16 (.Y(G314),.A(G1),.B(G5));
NAND2X1 NAND2_17 (.Y(G317),.A(G9),.B(G13));
NAND2X1 NAND2_18 (.Y(G320),.A(G2),.B(G6));
NAND2X1 NAND2_19 (.Y(G323),.A(G10),.B(G14));
NAND2X1 NAND2_20 (.Y(G326),.A(G3),.B(G7));
NAND2X1 NAND2_21 (.Y(G329),.A(G11),.B(G15));
NAND2X1 NAND2_22 (.Y(G332),.A(G4),.B(G8));
NAND2X1 NAND2_23 (.Y(G335),.A(G12),.B(G16));
NAND2X1 NAND2_24 (.Y(G338),.A(G17),.B(G21));
NAND2X1 NAND2_25 (.Y(G341),.A(G25),.B(G29));
NAND2X1 NAND2_26 (.Y(G344),.A(G18),.B(G22));
NAND2X1 NAND2_27 (.Y(G347),.A(G26),.B(G30));
NAND2X1 NAND2_28 (.Y(G350),.A(G19),.B(G23));
NAND2X1 NAND2_29 (.Y(G353),.A(G27),.B(G31));
NAND2X1 NAND2_30 (.Y(G356),.A(G20),.B(G24));
NAND2X1 NAND2_31 (.Y(G359),.A(G28),.B(G32));
NAND2X1 NAND2_32 (.Y(G362),.A(G1),.B(G266));
NAND2X1 NAND2_33 (.Y(G363),.A(G2),.B(G266));
NAND2X1 NAND2_34 (.Y(G364),.A(G3),.B(G269));
NAND2X1 NAND2_35 (.Y(G365),.A(G4),.B(G269));
NAND2X1 NAND2_36 (.Y(G366),.A(G5),.B(G272));
NAND2X1 NAND2_37 (.Y(G367),.A(G6),.B(G272));
NAND2X1 NAND2_38 (.Y(G368),.A(G7),.B(G275));
NAND2X1 NAND2_39 (.Y(G369),.A(G8),.B(G275));
NAND2X1 NAND2_40 (.Y(G370),.A(G9),.B(G278));
NAND2X1 NAND2_41 (.Y(G371),.A(G10),.B(G278));
NAND2X1 NAND2_42 (.Y(G372),.A(G11),.B(G281));
NAND2X1 NAND2_43 (.Y(G373),.A(G12),.B(G281));
NAND2X1 NAND2_44 (.Y(G374),.A(G13),.B(G284));
NAND2X1 NAND2_45 (.Y(G375),.A(G14),.B(G284));
NAND2X1 NAND2_46 (.Y(G376),.A(G15),.B(G287));
NAND2X1 NAND2_47 (.Y(G377),.A(G16),.B(G287));
NAND2X1 NAND2_48 (.Y(G378),.A(G17),.B(G290));
NAND2X1 NAND2_49 (.Y(G379),.A(G18),.B(G290));
NAND2X1 NAND2_50 (.Y(G380),.A(G19),.B(G293));
NAND2X1 NAND2_51 (.Y(G381),.A(G20),.B(G293));
NAND2X1 NAND2_52 (.Y(G382),.A(G21),.B(G296));
NAND2X1 NAND2_53 (.Y(G383),.A(G22),.B(G296));
NAND2X1 NAND2_54 (.Y(G384),.A(G23),.B(G299));
NAND2X1 NAND2_55 (.Y(G385),.A(G24),.B(G299));
NAND2X1 NAND2_56 (.Y(G386),.A(G25),.B(G302));
NAND2X1 NAND2_57 (.Y(G387),.A(G26),.B(G302));
NAND2X1 NAND2_58 (.Y(G388),.A(G27),.B(G305));
NAND2X1 NAND2_59 (.Y(G389),.A(G28),.B(G305));
NAND2X1 NAND2_60 (.Y(G390),.A(G29),.B(G308));
NAND2X1 NAND2_61 (.Y(G391),.A(G30),.B(G308));
NAND2X1 NAND2_62 (.Y(G392),.A(G31),.B(G311));
NAND2X1 NAND2_63 (.Y(G393),.A(G32),.B(G311));
NAND2X1 NAND2_64 (.Y(G394),.A(G1),.B(G314));
NAND2X1 NAND2_65 (.Y(G395),.A(G5),.B(G314));
NAND2X1 NAND2_66 (.Y(G396),.A(G9),.B(G317));
NAND2X1 NAND2_67 (.Y(G397),.A(G13),.B(G317));
NAND2X1 NAND2_68 (.Y(G398),.A(G2),.B(G320));
NAND2X1 NAND2_69 (.Y(G399),.A(G6),.B(G320));
NAND2X1 NAND2_70 (.Y(G400),.A(G10),.B(G323));
NAND2X1 NAND2_71 (.Y(G401),.A(G14),.B(G323));
NAND2X1 NAND2_72 (.Y(G402),.A(G3),.B(G326));
NAND2X1 NAND2_73 (.Y(G403),.A(G7),.B(G326));
NAND2X1 NAND2_74 (.Y(G404),.A(G11),.B(G329));
NAND2X1 NAND2_75 (.Y(G405),.A(G15),.B(G329));
NAND2X1 NAND2_76 (.Y(G406),.A(G4),.B(G332));
NAND2X1 NAND2_77 (.Y(G407),.A(G8),.B(G332));
NAND2X1 NAND2_78 (.Y(G408),.A(G12),.B(G335));
NAND2X1 NAND2_79 (.Y(G409),.A(G16),.B(G335));
NAND2X1 NAND2_80 (.Y(G410),.A(G17),.B(G338));
NAND2X1 NAND2_81 (.Y(G411),.A(G21),.B(G338));
NAND2X1 NAND2_82 (.Y(G412),.A(G25),.B(G341));
NAND2X1 NAND2_83 (.Y(G413),.A(G29),.B(G341));
NAND2X1 NAND2_84 (.Y(G414),.A(G18),.B(G344));
NAND2X1 NAND2_85 (.Y(G415),.A(G22),.B(G344));
NAND2X1 NAND2_86 (.Y(G416),.A(G26),.B(G347));
NAND2X1 NAND2_87 (.Y(G417),.A(G30),.B(G347));
NAND2X1 NAND2_88 (.Y(G418),.A(G19),.B(G350));
NAND2X1 NAND2_89 (.Y(G419),.A(G23),.B(G350));
NAND2X1 NAND2_90 (.Y(G420),.A(G27),.B(G353));
NAND2X1 NAND2_91 (.Y(G421),.A(G31),.B(G353));
NAND2X1 NAND2_92 (.Y(G422),.A(G20),.B(G356));
NAND2X1 NAND2_93 (.Y(G423),.A(G24),.B(G356));
NAND2X1 NAND2_94 (.Y(G424),.A(G28),.B(G359));
NAND2X1 NAND2_95 (.Y(G425),.A(G32),.B(G359));
NAND2X1 NAND2_96 (.Y(G426),.A(G362),.B(G363));
NAND2X1 NAND2_97 (.Y(G429),.A(G364),.B(G365));
NAND2X1 NAND2_98 (.Y(G432),.A(G366),.B(G367));
NAND2X1 NAND2_99 (.Y(G435),.A(G368),.B(G369));
NAND2X1 NAND2_100 (.Y(G438),.A(G370),.B(G371));
NAND2X1 NAND2_101 (.Y(G441),.A(G372),.B(G373));
NAND2X1 NAND2_102 (.Y(G444),.A(G374),.B(G375));
NAND2X1 NAND2_103 (.Y(G447),.A(G376),.B(G377));
NAND2X1 NAND2_104 (.Y(G450),.A(G378),.B(G379));
NAND2X1 NAND2_105 (.Y(G453),.A(G380),.B(G381));
NAND2X1 NAND2_106 (.Y(G456),.A(G382),.B(G383));
NAND2X1 NAND2_107 (.Y(G459),.A(G384),.B(G385));
NAND2X1 NAND2_108 (.Y(G462),.A(G386),.B(G387));
NAND2X1 NAND2_109 (.Y(G465),.A(G388),.B(G389));
NAND2X1 NAND2_110 (.Y(G468),.A(G390),.B(G391));
NAND2X1 NAND2_111 (.Y(G471),.A(G392),.B(G393));
NAND2X1 NAND2_112 (.Y(G474),.A(G394),.B(G395));
NAND2X1 NAND2_113 (.Y(G477),.A(G396),.B(G397));
NAND2X1 NAND2_114 (.Y(G480),.A(G398),.B(G399));
NAND2X1 NAND2_115 (.Y(G483),.A(G400),.B(G401));
NAND2X1 NAND2_116 (.Y(G486),.A(G402),.B(G403));
NAND2X1 NAND2_117 (.Y(G489),.A(G404),.B(G405));
NAND2X1 NAND2_118 (.Y(G492),.A(G406),.B(G407));
NAND2X1 NAND2_119 (.Y(G495),.A(G408),.B(G409));
NAND2X1 NAND2_120 (.Y(G498),.A(G410),.B(G411));
NAND2X1 NAND2_121 (.Y(G501),.A(G412),.B(G413));
NAND2X1 NAND2_122 (.Y(G504),.A(G414),.B(G415));
NAND2X1 NAND2_123 (.Y(G507),.A(G416),.B(G417));
NAND2X1 NAND2_124 (.Y(G510),.A(G418),.B(G419));
NAND2X1 NAND2_125 (.Y(G513),.A(G420),.B(G421));
NAND2X1 NAND2_126 (.Y(G516),.A(G422),.B(G423));
NAND2X1 NAND2_127 (.Y(G519),.A(G424),.B(G425));
NAND2X1 NAND2_128 (.Y(G522),.A(G426),.B(G429));
NAND2X1 NAND2_129 (.Y(G525),.A(G432),.B(G435));
NAND2X1 NAND2_130 (.Y(G528),.A(G438),.B(G441));
NAND2X1 NAND2_131 (.Y(G531),.A(G444),.B(G447));
NAND2X1 NAND2_132 (.Y(G534),.A(G450),.B(G453));
NAND2X1 NAND2_133 (.Y(G537),.A(G456),.B(G459));
NAND2X1 NAND2_134 (.Y(G540),.A(G462),.B(G465));
NAND2X1 NAND2_135 (.Y(G543),.A(G468),.B(G471));
NAND2X1 NAND2_136 (.Y(G546),.A(G474),.B(G477));
NAND2X1 NAND2_137 (.Y(G549),.A(G480),.B(G483));
NAND2X1 NAND2_138 (.Y(G552),.A(G486),.B(G489));
NAND2X1 NAND2_139 (.Y(G555),.A(G492),.B(G495));
NAND2X1 NAND2_140 (.Y(G558),.A(G498),.B(G501));
NAND2X1 NAND2_141 (.Y(G561),.A(G504),.B(G507));
NAND2X1 NAND2_142 (.Y(G564),.A(G510),.B(G513));
NAND2X1 NAND2_143 (.Y(G567),.A(G516),.B(G519));
NAND2X1 NAND2_144 (.Y(G570),.A(G426),.B(G522));
NAND2X1 NAND2_145 (.Y(G571),.A(G429),.B(G522));
NAND2X1 NAND2_146 (.Y(G572),.A(G432),.B(G525));
NAND2X1 NAND2_147 (.Y(G573),.A(G435),.B(G525));
NAND2X1 NAND2_148 (.Y(G574),.A(G438),.B(G528));
NAND2X1 NAND2_149 (.Y(G575),.A(G441),.B(G528));
NAND2X1 NAND2_150 (.Y(G576),.A(G444),.B(G531));
NAND2X1 NAND2_151 (.Y(G577),.A(G447),.B(G531));
NAND2X1 NAND2_152 (.Y(G578),.A(G450),.B(G534));
NAND2X1 NAND2_153 (.Y(G579),.A(G453),.B(G534));
NAND2X1 NAND2_154 (.Y(G580),.A(G456),.B(G537));
NAND2X1 NAND2_155 (.Y(G581),.A(G459),.B(G537));
NAND2X1 NAND2_156 (.Y(G582),.A(G462),.B(G540));
NAND2X1 NAND2_157 (.Y(G583),.A(G465),.B(G540));
NAND2X1 NAND2_158 (.Y(G584),.A(G468),.B(G543));
NAND2X1 NAND2_159 (.Y(G585),.A(G471),.B(G543));
NAND2X1 NAND2_160 (.Y(G586),.A(G474),.B(G546));
NAND2X1 NAND2_161 (.Y(G587),.A(G477),.B(G546));
NAND2X1 NAND2_162 (.Y(G588),.A(G480),.B(G549));
NAND2X1 NAND2_163 (.Y(G589),.A(G483),.B(G549));
NAND2X1 NAND2_164 (.Y(G590),.A(G486),.B(G552));
NAND2X1 NAND2_165 (.Y(G591),.A(G489),.B(G552));
NAND2X1 NAND2_166 (.Y(G592),.A(G492),.B(G555));
NAND2X1 NAND2_167 (.Y(G593),.A(G495),.B(G555));
NAND2X1 NAND2_168 (.Y(G594),.A(G498),.B(G558));
NAND2X1 NAND2_169 (.Y(G595),.A(G501),.B(G558));
NAND2X1 NAND2_170 (.Y(G596),.A(G504),.B(G561));
NAND2X1 NAND2_171 (.Y(G597),.A(G507),.B(G561));
NAND2X1 NAND2_172 (.Y(G598),.A(G510),.B(G564));
NAND2X1 NAND2_173 (.Y(G599),.A(G513),.B(G564));
NAND2X1 NAND2_174 (.Y(G600),.A(G516),.B(G567));
NAND2X1 NAND2_175 (.Y(G601),.A(G519),.B(G567));
NAND2X1 NAND2_176 (.Y(G602),.A(G570),.B(G571));
NAND2X1 NAND2_177 (.Y(G607),.A(G572),.B(G573));
NAND2X1 NAND2_178 (.Y(G612),.A(G574),.B(G575));
NAND2X1 NAND2_179 (.Y(G617),.A(G576),.B(G577));
NAND2X1 NAND2_180 (.Y(G622),.A(G578),.B(G579));
NAND2X1 NAND2_181 (.Y(G627),.A(G580),.B(G581));
NAND2X1 NAND2_182 (.Y(G632),.A(G582),.B(G583));
NAND2X1 NAND2_183 (.Y(G637),.A(G584),.B(G585));
NAND2X1 NAND2_184 (.Y(G642),.A(G586),.B(G587));
NAND2X1 NAND2_185 (.Y(G645),.A(G588),.B(G589));
NAND2X1 NAND2_186 (.Y(G648),.A(G590),.B(G591));
NAND2X1 NAND2_187 (.Y(G651),.A(G592),.B(G593));
NAND2X1 NAND2_188 (.Y(G654),.A(G594),.B(G595));
NAND2X1 NAND2_189 (.Y(G657),.A(G596),.B(G597));
NAND2X1 NAND2_190 (.Y(G660),.A(G598),.B(G599));
NAND2X1 NAND2_191 (.Y(G663),.A(G600),.B(G601));
NAND2X1 NAND2_192 (.Y(G666),.A(G602),.B(G607));
NAND2X1 NAND2_193 (.Y(G669),.A(G612),.B(G617));
NAND2X1 NAND2_194 (.Y(G672),.A(G602),.B(G612));
NAND2X1 NAND2_195 (.Y(G675),.A(G607),.B(G617));
NAND2X1 NAND2_196 (.Y(G678),.A(G622),.B(G627));
NAND2X1 NAND2_197 (.Y(G681),.A(G632),.B(G637));
NAND2X1 NAND2_198 (.Y(G684),.A(G622),.B(G632));
NAND2X1 NAND2_199 (.Y(G687),.A(G627),.B(G637));
NAND2X1 NAND2_200 (.Y(G690),.A(G602),.B(G666));
NAND2X1 NAND2_201 (.Y(G691),.A(G607),.B(G666));
NAND2X1 NAND2_202 (.Y(G692),.A(G612),.B(G669));
NAND2X1 NAND2_203 (.Y(G693),.A(G617),.B(G669));
NAND2X1 NAND2_204 (.Y(G694),.A(G602),.B(G672));
NAND2X1 NAND2_205 (.Y(G695),.A(G612),.B(G672));
NAND2X1 NAND2_206 (.Y(G696),.A(G607),.B(G675));
NAND2X1 NAND2_207 (.Y(G697),.A(G617),.B(G675));
NAND2X1 NAND2_208 (.Y(G698),.A(G622),.B(G678));
NAND2X1 NAND2_209 (.Y(G699),.A(G627),.B(G678));
NAND2X1 NAND2_210 (.Y(G700),.A(G632),.B(G681));
NAND2X1 NAND2_211 (.Y(G701),.A(G637),.B(G681));
NAND2X1 NAND2_212 (.Y(G702),.A(G622),.B(G684));
NAND2X1 NAND2_213 (.Y(G703),.A(G632),.B(G684));
NAND2X1 NAND2_214 (.Y(G704),.A(G627),.B(G687));
NAND2X1 NAND2_215 (.Y(G705),.A(G637),.B(G687));
NAND2X1 NAND2_216 (.Y(G706),.A(G690),.B(G691));
NAND2X1 NAND2_217 (.Y(G709),.A(G692),.B(G693));
NAND2X1 NAND2_218 (.Y(G712),.A(G694),.B(G695));
NAND2X1 NAND2_219 (.Y(G715),.A(G696),.B(G697));
NAND2X1 NAND2_220 (.Y(G718),.A(G698),.B(G699));
NAND2X1 NAND2_221 (.Y(G721),.A(G700),.B(G701));
NAND2X1 NAND2_222 (.Y(G724),.A(G702),.B(G703));
NAND2X1 NAND2_223 (.Y(G727),.A(G704),.B(G705));
NAND2X1 NAND2_224 (.Y(G730),.A(G242),.B(G718));
NAND2X1 NAND2_225 (.Y(G733),.A(G245),.B(G721));
NAND2X1 NAND2_226 (.Y(G736),.A(G248),.B(G724));
NAND2X1 NAND2_227 (.Y(G739),.A(G251),.B(G727));
NAND2X1 NAND2_228 (.Y(G742),.A(G254),.B(G706));
NAND2X1 NAND2_229 (.Y(G745),.A(G257),.B(G709));
NAND2X1 NAND2_230 (.Y(G748),.A(G260),.B(G712));
NAND2X1 NAND2_231 (.Y(G751),.A(G263),.B(G715));
NAND2X1 NAND2_232 (.Y(G754),.A(G242),.B(G730));
NAND2X1 NAND2_233 (.Y(G755),.A(G718),.B(G730));
NAND2X1 NAND2_234 (.Y(G756),.A(G245),.B(G733));
NAND2X1 NAND2_235 (.Y(G757),.A(G721),.B(G733));
NAND2X1 NAND2_236 (.Y(G758),.A(G248),.B(G736));
NAND2X1 NAND2_237 (.Y(G759),.A(G724),.B(G736));
NAND2X1 NAND2_238 (.Y(G760),.A(G251),.B(G739));
NAND2X1 NAND2_239 (.Y(G761),.A(G727),.B(G739));
NAND2X1 NAND2_240 (.Y(G762),.A(G254),.B(G742));
NAND2X1 NAND2_241 (.Y(G763),.A(G706),.B(G742));
NAND2X1 NAND2_242 (.Y(G764),.A(G257),.B(G745));
NAND2X1 NAND2_243 (.Y(G765),.A(G709),.B(G745));
NAND2X1 NAND2_244 (.Y(G766),.A(G260),.B(G748));
NAND2X1 NAND2_245 (.Y(G767),.A(G712),.B(G748));
NAND2X1 NAND2_246 (.Y(G768),.A(G263),.B(G751));
NAND2X1 NAND2_247 (.Y(G769),.A(G715),.B(G751));
NAND2X1 NAND2_248 (.Y(G770),.A(G754),.B(G755));
NAND2X1 NAND2_249 (.Y(G773),.A(G756),.B(G757));
NAND2X1 NAND2_250 (.Y(G776),.A(G758),.B(G759));
NAND2X1 NAND2_251 (.Y(G779),.A(G760),.B(G761));
NAND2X1 NAND2_252 (.Y(G782),.A(G762),.B(G763));
NAND2X1 NAND2_253 (.Y(G785),.A(G764),.B(G765));
NAND2X1 NAND2_254 (.Y(G788),.A(G766),.B(G767));
NAND2X1 NAND2_255 (.Y(G791),.A(G768),.B(G769));
NAND2X1 NAND2_256 (.Y(G794),.A(G642),.B(G770));
NAND2X1 NAND2_257 (.Y(G797),.A(G645),.B(G773));
NAND2X1 NAND2_258 (.Y(G800),.A(G648),.B(G776));
NAND2X1 NAND2_259 (.Y(G803),.A(G651),.B(G779));
NAND2X1 NAND2_260 (.Y(G806),.A(G654),.B(G782));
NAND2X1 NAND2_261 (.Y(G809),.A(G657),.B(G785));
NAND2X1 NAND2_262 (.Y(G812),.A(G660),.B(G788));
NAND2X1 NAND2_263 (.Y(G815),.A(G663),.B(G791));
NAND2X1 NAND2_264 (.Y(G818),.A(G642),.B(G794));
NAND2X1 NAND2_265 (.Y(G819),.A(G770),.B(G794));
NAND2X1 NAND2_266 (.Y(G820),.A(G645),.B(G797));
NAND2X1 NAND2_267 (.Y(G821),.A(G773),.B(G797));
NAND2X1 NAND2_268 (.Y(G822),.A(G648),.B(G800));
NAND2X1 NAND2_269 (.Y(G823),.A(G776),.B(G800));
NAND2X1 NAND2_270 (.Y(G824),.A(G651),.B(G803));
NAND2X1 NAND2_271 (.Y(G825),.A(G779),.B(G803));
NAND2X1 NAND2_272 (.Y(G826),.A(G654),.B(G806));
NAND2X1 NAND2_273 (.Y(G827),.A(G782),.B(G806));
NAND2X1 NAND2_274 (.Y(G828),.A(G657),.B(G809));
NAND2X1 NAND2_275 (.Y(G829),.A(G785),.B(G809));
NAND2X1 NAND2_276 (.Y(G830),.A(G660),.B(G812));
NAND2X1 NAND2_277 (.Y(G831),.A(G788),.B(G812));
NAND2X1 NAND2_278 (.Y(G832),.A(G663),.B(G815));
NAND2X1 NAND2_279 (.Y(G833),.A(G791),.B(G815));
NAND2X1 NAND2_280 (.Y(G834),.A(G818),.B(G819));
NAND2X1 NAND2_281 (.Y(G847),.A(G820),.B(G821));
NAND2X1 NAND2_282 (.Y(G860),.A(G822),.B(G823));
NAND2X1 NAND2_283 (.Y(G873),.A(G824),.B(G825));
NAND2X1 NAND2_284 (.Y(G886),.A(G828),.B(G829));
NAND2X1 NAND2_285 (.Y(G899),.A(G832),.B(G833));
NAND2X1 NAND2_286 (.Y(G912),.A(G830),.B(G831));
NAND2X1 NAND2_287 (.Y(G925),.A(G826),.B(G827));
INVX1 NOT_0 (.Y(G938),.A(G834));
INVX1 NOT_1 (.Y(G939),.A(G847));
INVX1 NOT_2 (.Y(G940),.A(G860));
INVX1 NOT_3 (.Y(G941),.A(G834));
INVX1 NOT_4 (.Y(G942),.A(G847));
INVX1 NOT_5 (.Y(G943),.A(G873));
INVX1 NOT_6 (.Y(G944),.A(G834));
INVX1 NOT_7 (.Y(G945),.A(G860));
INVX1 NOT_8 (.Y(G946),.A(G873));
INVX1 NOT_9 (.Y(G947),.A(G847));
INVX1 NOT_10 (.Y(G948),.A(G860));
INVX1 NOT_11 (.Y(G949),.A(G873));
INVX1 NOT_12 (.Y(G950),.A(G886));
INVX1 NOT_13 (.Y(G951),.A(G899));
INVX1 NOT_14 (.Y(G952),.A(G886));
INVX1 NOT_15 (.Y(G953),.A(G912));
INVX1 NOT_16 (.Y(G954),.A(G925));
INVX1 NOT_17 (.Y(G955),.A(G899));
INVX1 NOT_18 (.Y(G956),.A(G925));
INVX1 NOT_19 (.Y(G957),.A(G912));
INVX1 NOT_20 (.Y(G958),.A(G925));
INVX1 NOT_21 (.Y(G959),.A(G886));
INVX1 NOT_22 (.Y(G960),.A(G912));
INVX1 NOT_23 (.Y(G961),.A(G925));
INVX1 NOT_24 (.Y(G962),.A(G886));
INVX1 NOT_25 (.Y(G963),.A(G899));
INVX1 NOT_26 (.Y(G964),.A(G925));
INVX1 NOT_27 (.Y(G965),.A(G912));
INVX1 NOT_28 (.Y(G966),.A(G899));
INVX1 NOT_29 (.Y(G967),.A(G886));
INVX1 NOT_30 (.Y(G968),.A(G912));
INVX1 NOT_31 (.Y(G969),.A(G899));
INVX1 NOT_32 (.Y(G970),.A(G847));
INVX1 NOT_33 (.Y(G971),.A(G873));
INVX1 NOT_34 (.Y(G972),.A(G847));
INVX1 NOT_35 (.Y(G973),.A(G860));
INVX1 NOT_36 (.Y(G974),.A(G834));
INVX1 NOT_37 (.Y(G975),.A(G873));
INVX1 NOT_38 (.Y(G976),.A(G834));
INVX1 NOT_39 (.Y(G977),.A(G860));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(G940),.B(G873));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(G938),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(G978),.A(G939),.B(ttmp2));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(G860),.B(G943));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(G941),.B(ttmp4));
AND2X1 AND_tmp6 (.Y(G979),.A(G942),.B(ttmp5));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(G945),.B(G946));
AND2X1 AND_tmp8 (.Y(ttmp8),.A(G944),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(G980),.A(G847),.B(ttmp8));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(G948),.B(G949));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(G834),.B(ttmp10));
AND2X1 AND_tmp12 (.Y(G981),.A(G947),.B(ttmp11));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(G960),.B(G899));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(G958),.B(ttmp13));
AND2X1 AND_tmp15 (.Y(G982),.A(G959),.B(ttmp14));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(G912),.B(G963));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(G961),.B(ttmp16));
AND2X1 AND_tmp18 (.Y(G983),.A(G962),.B(ttmp17));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(G965),.B(G966));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(G964),.B(ttmp19));
AND2X1 AND_tmp21 (.Y(G984),.A(G886),.B(ttmp20));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(G968),.B(G969));
AND2X1 AND_tmp23 (.Y(ttmp23),.A(G925),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(G985),.A(G967),.B(ttmp23));
OR2X1 OR_tmp25 (.Y(ttmp25),.A(G980),.B(G981));
OR2X1 OR_tmp26 (.Y(ttmp26),.A(G978),.B(ttmp25));
OR2X1 OR_tmp27 (.Y(G986),.A(G979),.B(ttmp26));
OR2X1 OR_tmp28 (.Y(ttmp28),.A(G984),.B(G985));
OR2X1 OR_tmp29 (.Y(ttmp29),.A(G982),.B(ttmp28));
OR2X1 OR_tmp30 (.Y(G991),.A(G983),.B(ttmp29));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(G951),.B(G986));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(G925),.B(ttmp31));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(G950),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(G996),.A(G912),.B(ttmp33));
AND2X1 AND_tmp35 (.Y(ttmp35),.A(G899),.B(G986));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(G925),.B(ttmp35));
AND2X1 AND_tmp37 (.Y(ttmp37),.A(G952),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(G1001),.A(G953),.B(ttmp37));
AND2X1 AND_tmp39 (.Y(ttmp39),.A(G955),.B(G986));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(G954),.B(ttmp39));
AND2X1 AND_tmp41 (.Y(ttmp41),.A(G886),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(G1006),.A(G912),.B(ttmp41));
AND2X1 AND_tmp43 (.Y(ttmp43),.A(G899),.B(G986));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(G956),.B(ttmp43));
AND2X1 AND_tmp45 (.Y(ttmp45),.A(G886),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(G1011),.A(G957),.B(ttmp45));
AND2X1 AND_tmp47 (.Y(ttmp47),.A(G971),.B(G991));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(G834),.B(ttmp47));
AND2X1 AND_tmp49 (.Y(ttmp49),.A(G970),.B(ttmp48));
AND2X1 AND_tmp50 (.Y(G1016),.A(G860),.B(ttmp49));
AND2X1 AND_tmp51 (.Y(ttmp51),.A(G873),.B(G991));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(G834),.B(ttmp51));
AND2X1 AND_tmp53 (.Y(ttmp53),.A(G972),.B(ttmp52));
AND2X1 AND_tmp54 (.Y(G1021),.A(G973),.B(ttmp53));
AND2X1 AND_tmp55 (.Y(ttmp55),.A(G975),.B(G991));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(G974),.B(ttmp55));
AND2X1 AND_tmp57 (.Y(ttmp57),.A(G847),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(G1026),.A(G860),.B(ttmp57));
AND2X1 AND_tmp59 (.Y(ttmp59),.A(G873),.B(G991));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(G976),.B(ttmp59));
AND2X1 AND_tmp61 (.Y(ttmp61),.A(G847),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(G1031),.A(G977),.B(ttmp61));
AND2X1 AND2_8 (.Y(G1036),.A(G834),.B(G996));
AND2X1 AND2_9 (.Y(G1039),.A(G847),.B(G996));
AND2X1 AND2_10 (.Y(G1042),.A(G860),.B(G996));
AND2X1 AND2_11 (.Y(G1045),.A(G873),.B(G996));
AND2X1 AND2_12 (.Y(G1048),.A(G834),.B(G1001));
AND2X1 AND2_13 (.Y(G1051),.A(G847),.B(G1001));
AND2X1 AND2_14 (.Y(G1054),.A(G860),.B(G1001));
AND2X1 AND2_15 (.Y(G1057),.A(G873),.B(G1001));
AND2X1 AND2_16 (.Y(G1060),.A(G834),.B(G1006));
AND2X1 AND2_17 (.Y(G1063),.A(G847),.B(G1006));
AND2X1 AND2_18 (.Y(G1066),.A(G860),.B(G1006));
AND2X1 AND2_19 (.Y(G1069),.A(G873),.B(G1006));
AND2X1 AND2_20 (.Y(G1072),.A(G834),.B(G1011));
AND2X1 AND2_21 (.Y(G1075),.A(G847),.B(G1011));
AND2X1 AND2_22 (.Y(G1078),.A(G860),.B(G1011));
AND2X1 AND2_23 (.Y(G1081),.A(G873),.B(G1011));
AND2X1 AND2_24 (.Y(G1084),.A(G925),.B(G1016));
AND2X1 AND2_25 (.Y(G1087),.A(G886),.B(G1016));
AND2X1 AND2_26 (.Y(G1090),.A(G912),.B(G1016));
AND2X1 AND2_27 (.Y(G1093),.A(G899),.B(G1016));
AND2X1 AND2_28 (.Y(G1096),.A(G925),.B(G1021));
AND2X1 AND2_29 (.Y(G1099),.A(G886),.B(G1021));
AND2X1 AND2_30 (.Y(G1102),.A(G912),.B(G1021));
AND2X1 AND2_31 (.Y(G1105),.A(G899),.B(G1021));
AND2X1 AND2_32 (.Y(G1108),.A(G925),.B(G1026));
AND2X1 AND2_33 (.Y(G1111),.A(G886),.B(G1026));
AND2X1 AND2_34 (.Y(G1114),.A(G912),.B(G1026));
AND2X1 AND2_35 (.Y(G1117),.A(G899),.B(G1026));
AND2X1 AND2_36 (.Y(G1120),.A(G925),.B(G1031));
AND2X1 AND2_37 (.Y(G1123),.A(G886),.B(G1031));
AND2X1 AND2_38 (.Y(G1126),.A(G912),.B(G1031));
AND2X1 AND2_39 (.Y(G1129),.A(G899),.B(G1031));
NAND2X1 NAND2_288 (.Y(G1132),.A(G1),.B(G1036));
NAND2X1 NAND2_289 (.Y(G1135),.A(G2),.B(G1039));
NAND2X1 NAND2_290 (.Y(G1138),.A(G3),.B(G1042));
NAND2X1 NAND2_291 (.Y(G1141),.A(G4),.B(G1045));
NAND2X1 NAND2_292 (.Y(G1144),.A(G5),.B(G1048));
NAND2X1 NAND2_293 (.Y(G1147),.A(G6),.B(G1051));
NAND2X1 NAND2_294 (.Y(G1150),.A(G7),.B(G1054));
NAND2X1 NAND2_295 (.Y(G1153),.A(G8),.B(G1057));
NAND2X1 NAND2_296 (.Y(G1156),.A(G9),.B(G1060));
NAND2X1 NAND2_297 (.Y(G1159),.A(G10),.B(G1063));
NAND2X1 NAND2_298 (.Y(G1162),.A(G11),.B(G1066));
NAND2X1 NAND2_299 (.Y(G1165),.A(G12),.B(G1069));
NAND2X1 NAND2_300 (.Y(G1168),.A(G13),.B(G1072));
NAND2X1 NAND2_301 (.Y(G1171),.A(G14),.B(G1075));
NAND2X1 NAND2_302 (.Y(G1174),.A(G15),.B(G1078));
NAND2X1 NAND2_303 (.Y(G1177),.A(G16),.B(G1081));
NAND2X1 NAND2_304 (.Y(G1180),.A(G17),.B(G1084));
NAND2X1 NAND2_305 (.Y(G1183),.A(G18),.B(G1087));
NAND2X1 NAND2_306 (.Y(G1186),.A(G19),.B(G1090));
NAND2X1 NAND2_307 (.Y(G1189),.A(G20),.B(G1093));
NAND2X1 NAND2_308 (.Y(G1192),.A(G21),.B(G1096));
NAND2X1 NAND2_309 (.Y(G1195),.A(G22),.B(G1099));
NAND2X1 NAND2_310 (.Y(G1198),.A(G23),.B(G1102));
NAND2X1 NAND2_311 (.Y(G1201),.A(G24),.B(G1105));
NAND2X1 NAND2_312 (.Y(G1204),.A(G25),.B(G1108));
NAND2X1 NAND2_313 (.Y(G1207),.A(G26),.B(G1111));
NAND2X1 NAND2_314 (.Y(G1210),.A(G27),.B(G1114));
NAND2X1 NAND2_315 (.Y(G1213),.A(G28),.B(G1117));
NAND2X1 NAND2_316 (.Y(G1216),.A(G29),.B(G1120));
NAND2X1 NAND2_317 (.Y(G1219),.A(G30),.B(G1123));
NAND2X1 NAND2_318 (.Y(G1222),.A(G31),.B(G1126));
NAND2X1 NAND2_319 (.Y(G1225),.A(G32),.B(G1129));
NAND2X1 NAND2_320 (.Y(G1228),.A(G1),.B(G1132));
NAND2X1 NAND2_321 (.Y(G1229),.A(G1036),.B(G1132));
NAND2X1 NAND2_322 (.Y(G1230),.A(G2),.B(G1135));
NAND2X1 NAND2_323 (.Y(G1231),.A(G1039),.B(G1135));
NAND2X1 NAND2_324 (.Y(G1232),.A(G3),.B(G1138));
NAND2X1 NAND2_325 (.Y(G1233),.A(G1042),.B(G1138));
NAND2X1 NAND2_326 (.Y(G1234),.A(G4),.B(G1141));
NAND2X1 NAND2_327 (.Y(G1235),.A(G1045),.B(G1141));
NAND2X1 NAND2_328 (.Y(G1236),.A(G5),.B(G1144));
NAND2X1 NAND2_329 (.Y(G1237),.A(G1048),.B(G1144));
NAND2X1 NAND2_330 (.Y(G1238),.A(G6),.B(G1147));
NAND2X1 NAND2_331 (.Y(G1239),.A(G1051),.B(G1147));
NAND2X1 NAND2_332 (.Y(G1240),.A(G7),.B(G1150));
NAND2X1 NAND2_333 (.Y(G1241),.A(G1054),.B(G1150));
NAND2X1 NAND2_334 (.Y(G1242),.A(G8),.B(G1153));
NAND2X1 NAND2_335 (.Y(G1243),.A(G1057),.B(G1153));
NAND2X1 NAND2_336 (.Y(G1244),.A(G9),.B(G1156));
NAND2X1 NAND2_337 (.Y(G1245),.A(G1060),.B(G1156));
NAND2X1 NAND2_338 (.Y(G1246),.A(G10),.B(G1159));
NAND2X1 NAND2_339 (.Y(G1247),.A(G1063),.B(G1159));
NAND2X1 NAND2_340 (.Y(G1248),.A(G11),.B(G1162));
NAND2X1 NAND2_341 (.Y(G1249),.A(G1066),.B(G1162));
NAND2X1 NAND2_342 (.Y(G1250),.A(G12),.B(G1165));
NAND2X1 NAND2_343 (.Y(G1251),.A(G1069),.B(G1165));
NAND2X1 NAND2_344 (.Y(G1252),.A(G13),.B(G1168));
NAND2X1 NAND2_345 (.Y(G1253),.A(G1072),.B(G1168));
NAND2X1 NAND2_346 (.Y(G1254),.A(G14),.B(G1171));
NAND2X1 NAND2_347 (.Y(G1255),.A(G1075),.B(G1171));
NAND2X1 NAND2_348 (.Y(G1256),.A(G15),.B(G1174));
NAND2X1 NAND2_349 (.Y(G1257),.A(G1078),.B(G1174));
NAND2X1 NAND2_350 (.Y(G1258),.A(G16),.B(G1177));
NAND2X1 NAND2_351 (.Y(G1259),.A(G1081),.B(G1177));
NAND2X1 NAND2_352 (.Y(G1260),.A(G17),.B(G1180));
NAND2X1 NAND2_353 (.Y(G1261),.A(G1084),.B(G1180));
NAND2X1 NAND2_354 (.Y(G1262),.A(G18),.B(G1183));
NAND2X1 NAND2_355 (.Y(G1263),.A(G1087),.B(G1183));
NAND2X1 NAND2_356 (.Y(G1264),.A(G19),.B(G1186));
NAND2X1 NAND2_357 (.Y(G1265),.A(G1090),.B(G1186));
NAND2X1 NAND2_358 (.Y(G1266),.A(G20),.B(G1189));
NAND2X1 NAND2_359 (.Y(G1267),.A(G1093),.B(G1189));
NAND2X1 NAND2_360 (.Y(G1268),.A(G21),.B(G1192));
NAND2X1 NAND2_361 (.Y(G1269),.A(G1096),.B(G1192));
NAND2X1 NAND2_362 (.Y(G1270),.A(G22),.B(G1195));
NAND2X1 NAND2_363 (.Y(G1271),.A(G1099),.B(G1195));
NAND2X1 NAND2_364 (.Y(G1272),.A(G23),.B(G1198));
NAND2X1 NAND2_365 (.Y(G1273),.A(G1102),.B(G1198));
NAND2X1 NAND2_366 (.Y(G1274),.A(G24),.B(G1201));
NAND2X1 NAND2_367 (.Y(G1275),.A(G1105),.B(G1201));
NAND2X1 NAND2_368 (.Y(G1276),.A(G25),.B(G1204));
NAND2X1 NAND2_369 (.Y(G1277),.A(G1108),.B(G1204));
NAND2X1 NAND2_370 (.Y(G1278),.A(G26),.B(G1207));
NAND2X1 NAND2_371 (.Y(G1279),.A(G1111),.B(G1207));
NAND2X1 NAND2_372 (.Y(G1280),.A(G27),.B(G1210));
NAND2X1 NAND2_373 (.Y(G1281),.A(G1114),.B(G1210));
NAND2X1 NAND2_374 (.Y(G1282),.A(G28),.B(G1213));
NAND2X1 NAND2_375 (.Y(G1283),.A(G1117),.B(G1213));
NAND2X1 NAND2_376 (.Y(G1284),.A(G29),.B(G1216));
NAND2X1 NAND2_377 (.Y(G1285),.A(G1120),.B(G1216));
NAND2X1 NAND2_378 (.Y(G1286),.A(G30),.B(G1219));
NAND2X1 NAND2_379 (.Y(G1287),.A(G1123),.B(G1219));
NAND2X1 NAND2_380 (.Y(G1288),.A(G31),.B(G1222));
NAND2X1 NAND2_381 (.Y(G1289),.A(G1126),.B(G1222));
NAND2X1 NAND2_382 (.Y(G1290),.A(G32),.B(G1225));
NAND2X1 NAND2_383 (.Y(G1291),.A(G1129),.B(G1225));
NAND2X1 NAND2_384 (.Y(G1292),.A(G1228),.B(G1229));
NAND2X1 NAND2_385 (.Y(G1293),.A(G1230),.B(G1231));
NAND2X1 NAND2_386 (.Y(G1294),.A(G1232),.B(G1233));
NAND2X1 NAND2_387 (.Y(G1295),.A(G1234),.B(G1235));
NAND2X1 NAND2_388 (.Y(G1296),.A(G1236),.B(G1237));
NAND2X1 NAND2_389 (.Y(G1297),.A(G1238),.B(G1239));
NAND2X1 NAND2_390 (.Y(G1298),.A(G1240),.B(G1241));
NAND2X1 NAND2_391 (.Y(G1299),.A(G1242),.B(G1243));
NAND2X1 NAND2_392 (.Y(G1300),.A(G1244),.B(G1245));
NAND2X1 NAND2_393 (.Y(G1301),.A(G1246),.B(G1247));
NAND2X1 NAND2_394 (.Y(G1302),.A(G1248),.B(G1249));
NAND2X1 NAND2_395 (.Y(G1303),.A(G1250),.B(G1251));
NAND2X1 NAND2_396 (.Y(G1304),.A(G1252),.B(G1253));
NAND2X1 NAND2_397 (.Y(G1305),.A(G1254),.B(G1255));
NAND2X1 NAND2_398 (.Y(G1306),.A(G1256),.B(G1257));
NAND2X1 NAND2_399 (.Y(G1307),.A(G1258),.B(G1259));
NAND2X1 NAND2_400 (.Y(G1308),.A(G1260),.B(G1261));
NAND2X1 NAND2_401 (.Y(G1309),.A(G1262),.B(G1263));
NAND2X1 NAND2_402 (.Y(G1310),.A(G1264),.B(G1265));
NAND2X1 NAND2_403 (.Y(G1311),.A(G1266),.B(G1267));
NAND2X1 NAND2_404 (.Y(G1312),.A(G1268),.B(G1269));
NAND2X1 NAND2_405 (.Y(G1313),.A(G1270),.B(G1271));
NAND2X1 NAND2_406 (.Y(G1314),.A(G1272),.B(G1273));
NAND2X1 NAND2_407 (.Y(G1315),.A(G1274),.B(G1275));
NAND2X1 NAND2_408 (.Y(G1316),.A(G1276),.B(G1277));
NAND2X1 NAND2_409 (.Y(G1317),.A(G1278),.B(G1279));
NAND2X1 NAND2_410 (.Y(G1318),.A(G1280),.B(G1281));
NAND2X1 NAND2_411 (.Y(G1319),.A(G1282),.B(G1283));
NAND2X1 NAND2_412 (.Y(G1320),.A(G1284),.B(G1285));
NAND2X1 NAND2_413 (.Y(G1321),.A(G1286),.B(G1287));
NAND2X1 NAND2_414 (.Y(G1322),.A(G1288),.B(G1289));
NAND2X1 NAND2_415 (.Y(G1323),.A(G1290),.B(G1291));
INVX1 NOT_40 (.Y(G1324),.A(G1292));
INVX1 NOT_41 (.Y(G1325),.A(G1293));
INVX1 NOT_42 (.Y(G1326),.A(G1294));
INVX1 NOT_43 (.Y(G1327),.A(G1295));
INVX1 NOT_44 (.Y(G1328),.A(G1296));
INVX1 NOT_45 (.Y(G1329),.A(G1297));
INVX1 NOT_46 (.Y(G1330),.A(G1298));
INVX1 NOT_47 (.Y(G1331),.A(G1299));
INVX1 NOT_48 (.Y(G1332),.A(G1300));
INVX1 NOT_49 (.Y(G1333),.A(G1301));
INVX1 NOT_50 (.Y(G1334),.A(G1302));
INVX1 NOT_51 (.Y(G1335),.A(G1303));
INVX1 NOT_52 (.Y(G1336),.A(G1304));
INVX1 NOT_53 (.Y(G1337),.A(G1305));
INVX1 NOT_54 (.Y(G1338),.A(G1306));
INVX1 NOT_55 (.Y(G1339),.A(G1307));
INVX1 NOT_56 (.Y(G1340),.A(G1308));
INVX1 NOT_57 (.Y(G1341),.A(G1309));
INVX1 NOT_58 (.Y(G1342),.A(G1310));
INVX1 NOT_59 (.Y(G1343),.A(G1311));
INVX1 NOT_60 (.Y(G1344),.A(G1312));
INVX1 NOT_61 (.Y(G1345),.A(G1313));
INVX1 NOT_62 (.Y(G1346),.A(G1314));
INVX1 NOT_63 (.Y(G1347),.A(G1315));
INVX1 NOT_64 (.Y(G1348),.A(G1316));
INVX1 NOT_65 (.Y(G1349),.A(G1317));
INVX1 NOT_66 (.Y(G1350),.A(G1318));
INVX1 NOT_67 (.Y(G1351),.A(G1319));
INVX1 NOT_68 (.Y(G1352),.A(G1320));
INVX1 NOT_69 (.Y(G1353),.A(G1321));
INVX1 NOT_70 (.Y(G1354),.A(G1322));
INVX1 NOT_71 (.Y(G1355),.A(G1323));
endmodule 