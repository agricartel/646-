module c2670 (N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O);
input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I;
output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;
wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877;
BUFX1 BUFF1_1 (.Y(N398),.A(N219));
BUFX1 BUFF1_2 (.Y(N400),.A(N219));
BUFX1 BUFF1_3 (.Y(N401),.A(N219));
AND2X1 AND2_4 (.Y(N405),.A(N1),.B(N3));
INVX1 NOT1_5 (.Y(N408),.A(N230));
BUFX1 BUFF1_6 (.Y(N419),.A(N253));
BUFX1 BUFF1_7 (.Y(N420),.A(N253));
INVX1 NOT1_8 (.Y(N425),.A(N262));
BUFX1 BUFF1_9 (.Y(N456),.A(N290));
BUFX1 BUFF1_10 (.Y(N457),.A(N290));
BUFX1 BUFF1_11 (.Y(N458),.A(N290));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N301),.B(N297));
AND2X1 AND_tmp2 (.Y(ttmp2),.A(N309),.B(ttmp1));
AND2X1 AND_tmp3 (.Y(N485),.A(N305),.B(ttmp2));
INVX1 NOT1_13 (.Y(N486),.A(N405));
INVX1 NOT1_14 (.Y(N487),.A(N44));
INVX1 NOT1_15 (.Y(N488),.A(N132));
INVX1 NOT1_16 (.Y(N489),.A(N82));
INVX1 NOT1_17 (.Y(N490),.A(N96));
INVX1 NOT1_18 (.Y(N491),.A(N69));
INVX1 NOT1_19 (.Y(N492),.A(N120));
INVX1 NOT1_20 (.Y(N493),.A(N57));
INVX1 NOT1_21 (.Y(N494),.A(N108));
AND2X1 AND_tmp4 (.Y(ttmp4),.A(N15),.B(N237));
AND2X1 AND_tmp5 (.Y(N495),.A(N2),.B(ttmp4));
BUFX1 BUFF1_23 (.Y(N496),.A(N237));
AND2X1 AND2_24 (.Y(N499),.A(N37),.B(N37));
BUFX1 BUFF1_25 (.Y(N500),.A(N219));
BUFX1 BUFF1_26 (.Y(N503),.A(N8));
BUFX1 BUFF1_27 (.Y(N506),.A(N8));
BUFX1 BUFF1_28 (.Y(N509),.A(N227));
BUFX1 BUFF1_29 (.Y(N521),.A(N234));
INVX1 NOT1_30 (.Y(N533),.A(N241));
INVX1 NOT1_31 (.Y(N537),.A(N246));
AND2X1 AND2_32 (.Y(N543),.A(N11),.B(N246));
AND2X1 AND_tmp6 (.Y(ttmp6),.A(N96),.B(N44));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N132),.B(ttmp6));
AND2X1 AND_tmp8 (.Y(N544),.A(N82),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(N108),.B(N69));
AND2X1 AND_tmp10 (.Y(ttmp10),.A(N120),.B(ttmp9));
AND2X1 AND_tmp11 (.Y(N547),.A(N57),.B(ttmp10));
BUFX1 BUFF1_35 (.Y(N550),.A(N227));
BUFX1 BUFF1_36 (.Y(N562),.A(N234));
INVX1 NOT1_37 (.Y(N574),.A(N256));
INVX1 NOT1_38 (.Y(N578),.A(N259));
BUFX1 BUFF1_39 (.Y(N582),.A(N319));
BUFX1 BUFF1_40 (.Y(N594),.A(N322));
INVX1 NOT1_41 (.Y(N606),.A(N328));
INVX1 NOT1_42 (.Y(N607),.A(N331));
INVX1 NOT1_43 (.Y(N608),.A(N334));
INVX1 NOT1_44 (.Y(N609),.A(N337));
INVX1 NOT1_45 (.Y(N610),.A(N340));
INVX1 NOT1_46 (.Y(N611),.A(N343));
INVX1 NOT1_47 (.Y(N612),.A(N352));
BUFX1 BUFF1_48 (.Y(N613),.A(N319));
BUFX1 BUFF1_49 (.Y(N625),.A(N322));
BUFX1 BUFF1_50 (.Y(N637),.A(N16));
BUFX1 BUFF1_51 (.Y(N643),.A(N16));
INVX1 NOT1_52 (.Y(N650),.A(N355));
AND2X1 AND2_53 (.Y(N651),.A(N7),.B(N237));
INVX1 NOT1_54 (.Y(N655),.A(N263));
INVX1 NOT1_55 (.Y(N659),.A(N266));
INVX1 NOT1_56 (.Y(N663),.A(N269));
INVX1 NOT1_57 (.Y(N667),.A(N272));
INVX1 NOT1_58 (.Y(N671),.A(N275));
INVX1 NOT1_59 (.Y(N675),.A(N278));
INVX1 NOT1_60 (.Y(N679),.A(N281));
INVX1 NOT1_61 (.Y(N683),.A(N284));
INVX1 NOT1_62 (.Y(N687),.A(N287));
BUFX1 BUFF1_63 (.Y(N693),.A(N29));
BUFX1 BUFF1_64 (.Y(N699),.A(N29));
INVX1 NOT1_65 (.Y(N705),.A(N294));
INVX1 NOT1_66 (.Y(N711),.A(N297));
INVX1 NOT1_67 (.Y(N715),.A(N301));
INVX1 NOT1_68 (.Y(N719),.A(N305));
INVX1 NOT1_69 (.Y(N723),.A(N309));
INVX1 NOT1_70 (.Y(N727),.A(N313));
INVX1 NOT1_71 (.Y(N730),.A(N316));
INVX1 NOT1_72 (.Y(N733),.A(N346));
INVX1 NOT1_73 (.Y(N734),.A(N349));
BUFX1 BUFF1_74 (.Y(N735),.A(N259));
BUFX1 BUFF1_75 (.Y(N738),.A(N256));
BUFX1 BUFF1_76 (.Y(N741),.A(N263));
BUFX1 BUFF1_77 (.Y(N744),.A(N269));
BUFX1 BUFF1_78 (.Y(N747),.A(N266));
BUFX1 BUFF1_79 (.Y(N750),.A(N275));
BUFX1 BUFF1_80 (.Y(N753),.A(N272));
BUFX1 BUFF1_81 (.Y(N756),.A(N281));
BUFX1 BUFF1_82 (.Y(N759),.A(N278));
BUFX1 BUFF1_83 (.Y(N762),.A(N287));
BUFX1 BUFF1_84 (.Y(N765),.A(N284));
BUFX1 BUFF1_85 (.Y(N768),.A(N294));
BUFX1 BUFF1_86 (.Y(N771),.A(N301));
BUFX1 BUFF1_87 (.Y(N774),.A(N297));
BUFX1 BUFF1_88 (.Y(N777),.A(N309));
BUFX1 BUFF1_89 (.Y(N780),.A(N305));
BUFX1 BUFF1_90 (.Y(N783),.A(N316));
BUFX1 BUFF1_91 (.Y(N786),.A(N313));
INVX1 NOT1_92 (.Y(N792),.A(N485));
INVX1 NOT1_93 (.Y(N799),.A(N495));
INVX1 NOT1_94 (.Y(N800),.A(N499));
BUFX1 BUFF1_95 (.Y(N805),.A(N500));
NAND2X1 NAND2_96 (.Y(N900),.A(N331),.B(N606));
NAND2X1 NAND2_97 (.Y(N901),.A(N328),.B(N607));
NAND2X1 NAND2_98 (.Y(N902),.A(N337),.B(N608));
NAND2X1 NAND2_99 (.Y(N903),.A(N334),.B(N609));
NAND2X1 NAND2_100 (.Y(N904),.A(N343),.B(N610));
NAND2X1 NAND2_101 (.Y(N905),.A(N340),.B(N611));
NAND2X1 NAND2_102 (.Y(N998),.A(N349),.B(N733));
NAND2X1 NAND2_103 (.Y(N999),.A(N346),.B(N734));
AND2X1 AND2_104 (.Y(N1026),.A(N94),.B(N500));
AND2X1 AND2_105 (.Y(N1027),.A(N325),.B(N651));
INVX1 NOT1_106 (.Y(N1028),.A(N651));
NAND2X1 NAND2_107 (.Y(N1029),.A(N231),.B(N651));
INVX1 NOT1_108 (.Y(N1032),.A(N544));
INVX1 NOT1_109 (.Y(N1033),.A(N547));
AND2X1 AND2_110 (.Y(N1034),.A(N547),.B(N544));
BUFX1 BUFF1_111 (.Y(N1037),.A(N503));
INVX1 NOT1_112 (.Y(N1042),.A(N509));
INVX1 NOT1_113 (.Y(N1053),.A(N521));
AND2X1 AND_tmp12 (.Y(ttmp12),.A(N509),.B(N521));
AND2X1 AND_tmp13 (.Y(N1064),.A(N80),.B(ttmp12));
AND2X1 AND_tmp14 (.Y(ttmp14),.A(N509),.B(N521));
AND2X1 AND_tmp15 (.Y(N1065),.A(N68),.B(ttmp14));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(N509),.B(N521));
AND2X1 AND_tmp17 (.Y(N1066),.A(N79),.B(ttmp16));
AND2X1 AND_tmp18 (.Y(ttmp18),.A(N509),.B(N521));
AND2X1 AND_tmp19 (.Y(N1067),.A(N78),.B(ttmp18));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(N509),.B(N521));
AND2X1 AND_tmp21 (.Y(N1068),.A(N77),.B(ttmp20));
AND2X1 AND2_119 (.Y(N1069),.A(N11),.B(N537));
BUFX1 BUFF1_120 (.Y(N1070),.A(N503));
INVX1 NOT1_121 (.Y(N1075),.A(N550));
INVX1 NOT1_122 (.Y(N1086),.A(N562));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N550),.B(N562));
AND2X1 AND_tmp23 (.Y(N1097),.A(N76),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N550),.B(N562));
AND2X1 AND_tmp25 (.Y(N1098),.A(N75),.B(ttmp24));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(N550),.B(N562));
AND2X1 AND_tmp27 (.Y(N1099),.A(N74),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(ttmp28),.A(N550),.B(N562));
AND2X1 AND_tmp29 (.Y(N1100),.A(N73),.B(ttmp28));
AND2X1 AND_tmp30 (.Y(ttmp30),.A(N550),.B(N562));
AND2X1 AND_tmp31 (.Y(N1101),.A(N72),.B(ttmp30));
INVX1 NOT1_128 (.Y(N1102),.A(N582));
INVX1 NOT1_129 (.Y(N1113),.A(N594));
AND2X1 AND_tmp32 (.Y(ttmp32),.A(N582),.B(N594));
AND2X1 AND_tmp33 (.Y(N1124),.A(N114),.B(ttmp32));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N582),.B(N594));
AND2X1 AND_tmp35 (.Y(N1125),.A(N113),.B(ttmp34));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N582),.B(N594));
AND2X1 AND_tmp37 (.Y(N1126),.A(N112),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N582),.B(N594));
AND2X1 AND_tmp39 (.Y(N1127),.A(N111),.B(ttmp38));
AND2X1 AND2_134 (.Y(N1128),.A(N582),.B(N594));
NAND2X1 NAND2_135 (.Y(N1129),.A(N900),.B(N901));
NAND2X1 NAND2_136 (.Y(N1133),.A(N902),.B(N903));
NAND2X1 NAND2_137 (.Y(N1137),.A(N904),.B(N905));
INVX1 NOT1_138 (.Y(N1140),.A(N741));
NAND2X1 NAND2_139 (.Y(N1141),.A(N741),.B(N612));
INVX1 NOT1_140 (.Y(N1142),.A(N744));
INVX1 NOT1_141 (.Y(N1143),.A(N747));
INVX1 NOT1_142 (.Y(N1144),.A(N750));
INVX1 NOT1_143 (.Y(N1145),.A(N753));
INVX1 NOT1_144 (.Y(N1146),.A(N613));
INVX1 NOT1_145 (.Y(N1157),.A(N625));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N613),.B(N625));
AND2X1 AND_tmp41 (.Y(N1168),.A(N118),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(N613),.B(N625));
AND2X1 AND_tmp43 (.Y(N1169),.A(N107),.B(ttmp42));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N613),.B(N625));
AND2X1 AND_tmp45 (.Y(N1170),.A(N117),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(N613),.B(N625));
AND2X1 AND_tmp47 (.Y(N1171),.A(N116),.B(ttmp46));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(N613),.B(N625));
AND2X1 AND_tmp49 (.Y(N1172),.A(N115),.B(ttmp48));
INVX1 NOT1_151 (.Y(N1173),.A(N637));
INVX1 NOT1_152 (.Y(N1178),.A(N643));
INVX1 NOT1_153 (.Y(N1184),.A(N768));
NAND2X1 NAND2_154 (.Y(N1185),.A(N768),.B(N650));
INVX1 NOT1_155 (.Y(N1186),.A(N771));
INVX1 NOT1_156 (.Y(N1187),.A(N774));
INVX1 NOT1_157 (.Y(N1188),.A(N777));
INVX1 NOT1_158 (.Y(N1189),.A(N780));
BUFX1 BUFF1_159 (.Y(N1190),.A(N506));
BUFX1 BUFF1_160 (.Y(N1195),.A(N506));
INVX1 NOT1_161 (.Y(N1200),.A(N693));
INVX1 NOT1_162 (.Y(N1205),.A(N699));
INVX1 NOT1_163 (.Y(N1210),.A(N735));
INVX1 NOT1_164 (.Y(N1211),.A(N738));
INVX1 NOT1_165 (.Y(N1212),.A(N756));
INVX1 NOT1_166 (.Y(N1213),.A(N759));
INVX1 NOT1_167 (.Y(N1214),.A(N762));
INVX1 NOT1_168 (.Y(N1215),.A(N765));
NAND2X1 NAND2_169 (.Y(N1216),.A(N998),.B(N999));
BUFX1 BUFF1_170 (.Y(N1219),.A(N574));
BUFX1 BUFF1_171 (.Y(N1222),.A(N578));
BUFX1 BUFF1_172 (.Y(N1225),.A(N655));
BUFX1 BUFF1_173 (.Y(N1228),.A(N659));
BUFX1 BUFF1_174 (.Y(N1231),.A(N663));
BUFX1 BUFF1_175 (.Y(N1234),.A(N667));
BUFX1 BUFF1_176 (.Y(N1237),.A(N671));
BUFX1 BUFF1_177 (.Y(N1240),.A(N675));
BUFX1 BUFF1_178 (.Y(N1243),.A(N679));
BUFX1 BUFF1_179 (.Y(N1246),.A(N683));
INVX1 NOT1_180 (.Y(N1249),.A(N783));
INVX1 NOT1_181 (.Y(N1250),.A(N786));
BUFX1 BUFF1_182 (.Y(N1251),.A(N687));
BUFX1 BUFF1_183 (.Y(N1254),.A(N705));
BUFX1 BUFF1_184 (.Y(N1257),.A(N711));
BUFX1 BUFF1_185 (.Y(N1260),.A(N715));
BUFX1 BUFF1_186 (.Y(N1263),.A(N719));
BUFX1 BUFF1_187 (.Y(N1266),.A(N723));
INVX1 NOT1_188 (.Y(N1269),.A(N1027));
AND2X1 AND2_189 (.Y(N1275),.A(N325),.B(N1032));
AND2X1 AND2_190 (.Y(N1276),.A(N231),.B(N1033));
BUFX1 BUFF1_191 (.Y(N1277),.A(N1034));
OR2X1 OR2_192 (.Y(N1302),.A(N1069),.B(N543));
NAND2X1 NAND2_193 (.Y(N1351),.A(N352),.B(N1140));
NAND2X1 NAND2_194 (.Y(N1352),.A(N747),.B(N1142));
NAND2X1 NAND2_195 (.Y(N1353),.A(N744),.B(N1143));
NAND2X1 NAND2_196 (.Y(N1354),.A(N753),.B(N1144));
NAND2X1 NAND2_197 (.Y(N1355),.A(N750),.B(N1145));
NAND2X1 NAND2_198 (.Y(N1395),.A(N355),.B(N1184));
NAND2X1 NAND2_199 (.Y(N1396),.A(N774),.B(N1186));
NAND2X1 NAND2_200 (.Y(N1397),.A(N771),.B(N1187));
NAND2X1 NAND2_201 (.Y(N1398),.A(N780),.B(N1188));
NAND2X1 NAND2_202 (.Y(N1399),.A(N777),.B(N1189));
NAND2X1 NAND2_203 (.Y(N1422),.A(N738),.B(N1210));
NAND2X1 NAND2_204 (.Y(N1423),.A(N735),.B(N1211));
NAND2X1 NAND2_205 (.Y(N1424),.A(N759),.B(N1212));
NAND2X1 NAND2_206 (.Y(N1425),.A(N756),.B(N1213));
NAND2X1 NAND2_207 (.Y(N1426),.A(N765),.B(N1214));
NAND2X1 NAND2_208 (.Y(N1427),.A(N762),.B(N1215));
NAND2X1 NAND2_209 (.Y(N1440),.A(N786),.B(N1249));
NAND2X1 NAND2_210 (.Y(N1441),.A(N783),.B(N1250));
INVX1 NOT1_211 (.Y(N1448),.A(N1034));
INVX1 NOT1_212 (.Y(N1449),.A(N1275));
INVX1 NOT1_213 (.Y(N1450),.A(N1276));
AND2X1 AND_tmp50 (.Y(ttmp50),.A(N1042),.B(N1053));
AND2X1 AND_tmp51 (.Y(N1451),.A(N93),.B(ttmp50));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(N509),.B(N1053));
AND2X1 AND_tmp53 (.Y(N1452),.A(N55),.B(ttmp52));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(N1042),.B(N521));
AND2X1 AND_tmp55 (.Y(N1453),.A(N67),.B(ttmp54));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(N1042),.B(N1053));
AND2X1 AND_tmp57 (.Y(N1454),.A(N81),.B(ttmp56));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(N509),.B(N1053));
AND2X1 AND_tmp59 (.Y(N1455),.A(N43),.B(ttmp58));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N1042),.B(N521));
AND2X1 AND_tmp61 (.Y(N1456),.A(N56),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N1042),.B(N1053));
AND2X1 AND_tmp63 (.Y(N1457),.A(N92),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(ttmp64),.A(N509),.B(N1053));
AND2X1 AND_tmp65 (.Y(N1458),.A(N54),.B(ttmp64));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(N1042),.B(N521));
AND2X1 AND_tmp67 (.Y(N1459),.A(N66),.B(ttmp66));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N1042),.B(N1053));
AND2X1 AND_tmp69 (.Y(N1460),.A(N91),.B(ttmp68));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N509),.B(N1053));
AND2X1 AND_tmp71 (.Y(N1461),.A(N53),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(ttmp72),.A(N1042),.B(N521));
AND2X1 AND_tmp73 (.Y(N1462),.A(N65),.B(ttmp72));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N1042),.B(N1053));
AND2X1 AND_tmp75 (.Y(N1463),.A(N90),.B(ttmp74));
AND2X1 AND_tmp76 (.Y(ttmp76),.A(N509),.B(N1053));
AND2X1 AND_tmp77 (.Y(N1464),.A(N52),.B(ttmp76));
AND2X1 AND_tmp78 (.Y(ttmp78),.A(N1042),.B(N521));
AND2X1 AND_tmp79 (.Y(N1465),.A(N64),.B(ttmp78));
AND2X1 AND_tmp80 (.Y(ttmp80),.A(N1075),.B(N1086));
AND2X1 AND_tmp81 (.Y(N1466),.A(N89),.B(ttmp80));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(N550),.B(N1086));
AND2X1 AND_tmp83 (.Y(N1467),.A(N51),.B(ttmp82));
AND2X1 AND_tmp84 (.Y(ttmp84),.A(N1075),.B(N562));
AND2X1 AND_tmp85 (.Y(N1468),.A(N63),.B(ttmp84));
AND2X1 AND_tmp86 (.Y(ttmp86),.A(N1075),.B(N1086));
AND2X1 AND_tmp87 (.Y(N1469),.A(N88),.B(ttmp86));
AND2X1 AND_tmp88 (.Y(ttmp88),.A(N550),.B(N1086));
AND2X1 AND_tmp89 (.Y(N1470),.A(N50),.B(ttmp88));
AND2X1 AND_tmp90 (.Y(ttmp90),.A(N1075),.B(N562));
AND2X1 AND_tmp91 (.Y(N1471),.A(N62),.B(ttmp90));
AND2X1 AND_tmp92 (.Y(ttmp92),.A(N1075),.B(N1086));
AND2X1 AND_tmp93 (.Y(N1472),.A(N87),.B(ttmp92));
AND2X1 AND_tmp94 (.Y(ttmp94),.A(N550),.B(N1086));
AND2X1 AND_tmp95 (.Y(N1473),.A(N49),.B(ttmp94));
AND2X1 AND2_237 (.Y(N1474),.A(N1075),.B(N562));
AND2X1 AND_tmp96 (.Y(ttmp96),.A(N1075),.B(N1086));
AND2X1 AND_tmp97 (.Y(N1475),.A(N86),.B(ttmp96));
AND2X1 AND_tmp98 (.Y(ttmp98),.A(N550),.B(N1086));
AND2X1 AND_tmp99 (.Y(N1476),.A(N48),.B(ttmp98));
AND2X1 AND_tmp100 (.Y(ttmp100),.A(N1075),.B(N562));
AND2X1 AND_tmp101 (.Y(N1477),.A(N61),.B(ttmp100));
AND2X1 AND_tmp102 (.Y(ttmp102),.A(N1075),.B(N1086));
AND2X1 AND_tmp103 (.Y(N1478),.A(N85),.B(ttmp102));
AND2X1 AND_tmp104 (.Y(ttmp104),.A(N550),.B(N1086));
AND2X1 AND_tmp105 (.Y(N1479),.A(N47),.B(ttmp104));
AND2X1 AND_tmp106 (.Y(ttmp106),.A(N1075),.B(N562));
AND2X1 AND_tmp107 (.Y(N1480),.A(N60),.B(ttmp106));
AND2X1 AND_tmp108 (.Y(ttmp108),.A(N1102),.B(N1113));
AND2X1 AND_tmp109 (.Y(N1481),.A(N138),.B(ttmp108));
AND2X1 AND_tmp110 (.Y(ttmp110),.A(N582),.B(N1113));
AND2X1 AND_tmp111 (.Y(N1482),.A(N102),.B(ttmp110));
AND2X1 AND_tmp112 (.Y(ttmp112),.A(N1102),.B(N594));
AND2X1 AND_tmp113 (.Y(N1483),.A(N126),.B(ttmp112));
AND2X1 AND_tmp114 (.Y(ttmp114),.A(N1102),.B(N1113));
AND2X1 AND_tmp115 (.Y(N1484),.A(N137),.B(ttmp114));
AND2X1 AND_tmp116 (.Y(ttmp116),.A(N582),.B(N1113));
AND2X1 AND_tmp117 (.Y(N1485),.A(N101),.B(ttmp116));
AND2X1 AND_tmp118 (.Y(ttmp118),.A(N1102),.B(N594));
AND2X1 AND_tmp119 (.Y(N1486),.A(N125),.B(ttmp118));
AND2X1 AND_tmp120 (.Y(ttmp120),.A(N1102),.B(N1113));
AND2X1 AND_tmp121 (.Y(N1487),.A(N136),.B(ttmp120));
AND2X1 AND_tmp122 (.Y(ttmp122),.A(N582),.B(N1113));
AND2X1 AND_tmp123 (.Y(N1488),.A(N100),.B(ttmp122));
AND2X1 AND_tmp124 (.Y(ttmp124),.A(N1102),.B(N594));
AND2X1 AND_tmp125 (.Y(N1489),.A(N124),.B(ttmp124));
AND2X1 AND_tmp126 (.Y(ttmp126),.A(N1102),.B(N1113));
AND2X1 AND_tmp127 (.Y(N1490),.A(N135),.B(ttmp126));
AND2X1 AND_tmp128 (.Y(ttmp128),.A(N582),.B(N1113));
AND2X1 AND_tmp129 (.Y(N1491),.A(N99),.B(ttmp128));
AND2X1 AND_tmp130 (.Y(ttmp130),.A(N1102),.B(N594));
AND2X1 AND_tmp131 (.Y(N1492),.A(N123),.B(ttmp130));
AND2X1 AND2_256 (.Y(N1493),.A(N1102),.B(N1113));
AND2X1 AND2_257 (.Y(N1494),.A(N582),.B(N1113));
AND2X1 AND2_258 (.Y(N1495),.A(N1102),.B(N594));
INVX1 NOT1_259 (.Y(N1496),.A(N1129));
INVX1 NOT1_260 (.Y(N1499),.A(N1133));
NAND2X1 NAND2_261 (.Y(N1502),.A(N1351),.B(N1141));
NAND2X1 NAND2_262 (.Y(N1506),.A(N1352),.B(N1353));
NAND2X1 NAND2_263 (.Y(N1510),.A(N1354),.B(N1355));
BUFX1 BUFF1_264 (.Y(N1513),.A(N1137));
BUFX1 BUFF1_265 (.Y(N1516),.A(N1137));
INVX1 NOT1_266 (.Y(N1519),.A(N1219));
INVX1 NOT1_267 (.Y(N1520),.A(N1222));
INVX1 NOT1_268 (.Y(N1521),.A(N1225));
INVX1 NOT1_269 (.Y(N1522),.A(N1228));
INVX1 NOT1_270 (.Y(N1523),.A(N1231));
INVX1 NOT1_271 (.Y(N1524),.A(N1234));
INVX1 NOT1_272 (.Y(N1525),.A(N1237));
INVX1 NOT1_273 (.Y(N1526),.A(N1240));
INVX1 NOT1_274 (.Y(N1527),.A(N1243));
INVX1 NOT1_275 (.Y(N1528),.A(N1246));
AND2X1 AND_tmp132 (.Y(ttmp132),.A(N1146),.B(N1157));
AND2X1 AND_tmp133 (.Y(N1529),.A(N142),.B(ttmp132));
AND2X1 AND_tmp134 (.Y(ttmp134),.A(N613),.B(N1157));
AND2X1 AND_tmp135 (.Y(N1530),.A(N106),.B(ttmp134));
AND2X1 AND_tmp136 (.Y(ttmp136),.A(N1146),.B(N625));
AND2X1 AND_tmp137 (.Y(N1531),.A(N130),.B(ttmp136));
AND2X1 AND_tmp138 (.Y(ttmp138),.A(N1146),.B(N1157));
AND2X1 AND_tmp139 (.Y(N1532),.A(N131),.B(ttmp138));
AND2X1 AND_tmp140 (.Y(ttmp140),.A(N613),.B(N1157));
AND2X1 AND_tmp141 (.Y(N1533),.A(N95),.B(ttmp140));
AND2X1 AND_tmp142 (.Y(ttmp142),.A(N1146),.B(N625));
AND2X1 AND_tmp143 (.Y(N1534),.A(N119),.B(ttmp142));
AND2X1 AND_tmp144 (.Y(ttmp144),.A(N1146),.B(N1157));
AND2X1 AND_tmp145 (.Y(N1535),.A(N141),.B(ttmp144));
AND2X1 AND_tmp146 (.Y(ttmp146),.A(N613),.B(N1157));
AND2X1 AND_tmp147 (.Y(N1536),.A(N105),.B(ttmp146));
AND2X1 AND_tmp148 (.Y(ttmp148),.A(N1146),.B(N625));
AND2X1 AND_tmp149 (.Y(N1537),.A(N129),.B(ttmp148));
AND2X1 AND_tmp150 (.Y(ttmp150),.A(N1146),.B(N1157));
AND2X1 AND_tmp151 (.Y(N1538),.A(N140),.B(ttmp150));
AND2X1 AND_tmp152 (.Y(ttmp152),.A(N613),.B(N1157));
AND2X1 AND_tmp153 (.Y(N1539),.A(N104),.B(ttmp152));
AND2X1 AND_tmp154 (.Y(ttmp154),.A(N1146),.B(N625));
AND2X1 AND_tmp155 (.Y(N1540),.A(N128),.B(ttmp154));
AND2X1 AND_tmp156 (.Y(ttmp156),.A(N1146),.B(N1157));
AND2X1 AND_tmp157 (.Y(N1541),.A(N139),.B(ttmp156));
AND2X1 AND_tmp158 (.Y(ttmp158),.A(N613),.B(N1157));
AND2X1 AND_tmp159 (.Y(N1542),.A(N103),.B(ttmp158));
AND2X1 AND_tmp160 (.Y(ttmp160),.A(N1146),.B(N625));
AND2X1 AND_tmp161 (.Y(N1543),.A(N127),.B(ttmp160));
AND2X1 AND2_291 (.Y(N1544),.A(N19),.B(N1173));
AND2X1 AND2_292 (.Y(N1545),.A(N4),.B(N1173));
AND2X1 AND2_293 (.Y(N1546),.A(N20),.B(N1173));
AND2X1 AND2_294 (.Y(N1547),.A(N5),.B(N1173));
AND2X1 AND2_295 (.Y(N1548),.A(N21),.B(N1178));
AND2X1 AND2_296 (.Y(N1549),.A(N22),.B(N1178));
AND2X1 AND2_297 (.Y(N1550),.A(N23),.B(N1178));
AND2X1 AND2_298 (.Y(N1551),.A(N6),.B(N1178));
AND2X1 AND2_299 (.Y(N1552),.A(N24),.B(N1178));
NAND2X1 NAND2_300 (.Y(N1553),.A(N1395),.B(N1185));
NAND2X1 NAND2_301 (.Y(N1557),.A(N1396),.B(N1397));
NAND2X1 NAND2_302 (.Y(N1561),.A(N1398),.B(N1399));
AND2X1 AND2_303 (.Y(N1564),.A(N25),.B(N1200));
AND2X1 AND2_304 (.Y(N1565),.A(N32),.B(N1200));
AND2X1 AND2_305 (.Y(N1566),.A(N26),.B(N1200));
AND2X1 AND2_306 (.Y(N1567),.A(N33),.B(N1200));
AND2X1 AND2_307 (.Y(N1568),.A(N27),.B(N1205));
AND2X1 AND2_308 (.Y(N1569),.A(N34),.B(N1205));
AND2X1 AND2_309 (.Y(N1570),.A(N35),.B(N1205));
AND2X1 AND2_310 (.Y(N1571),.A(N28),.B(N1205));
INVX1 NOT1_311 (.Y(N1572),.A(N1251));
INVX1 NOT1_312 (.Y(N1573),.A(N1254));
INVX1 NOT1_313 (.Y(N1574),.A(N1257));
INVX1 NOT1_314 (.Y(N1575),.A(N1260));
INVX1 NOT1_315 (.Y(N1576),.A(N1263));
INVX1 NOT1_316 (.Y(N1577),.A(N1266));
NAND2X1 NAND2_317 (.Y(N1578),.A(N1422),.B(N1423));
INVX1 NOT1_318 (.Y(N1581),.A(N1216));
NAND2X1 NAND2_319 (.Y(N1582),.A(N1426),.B(N1427));
NAND2X1 NAND2_320 (.Y(N1585),.A(N1424),.B(N1425));
NAND2X1 NAND2_321 (.Y(N1588),.A(N1440),.B(N1441));
AND2X1 AND2_322 (.Y(N1591),.A(N1449),.B(N1450));
OR2X1 OR_tmp162 (.Y(ttmp162),.A(N1453),.B(N1064));
OR2X1 OR_tmp163 (.Y(ttmp163),.A(N1451),.B(ttmp162));
OR2X1 OR_tmp164 (.Y(N1596),.A(N1452),.B(ttmp163));
OR2X1 OR_tmp165 (.Y(ttmp165),.A(N1456),.B(N1065));
OR2X1 OR_tmp166 (.Y(ttmp166),.A(N1454),.B(ttmp165));
OR2X1 OR_tmp167 (.Y(N1600),.A(N1455),.B(ttmp166));
OR2X1 OR_tmp168 (.Y(ttmp168),.A(N1459),.B(N1066));
OR2X1 OR_tmp169 (.Y(ttmp169),.A(N1457),.B(ttmp168));
OR2X1 OR_tmp170 (.Y(N1606),.A(N1458),.B(ttmp169));
OR2X1 OR_tmp171 (.Y(ttmp171),.A(N1462),.B(N1067));
OR2X1 OR_tmp172 (.Y(ttmp172),.A(N1460),.B(ttmp171));
OR2X1 OR_tmp173 (.Y(N1612),.A(N1461),.B(ttmp172));
OR2X1 OR_tmp174 (.Y(ttmp174),.A(N1465),.B(N1068));
OR2X1 OR_tmp175 (.Y(ttmp175),.A(N1463),.B(ttmp174));
OR2X1 OR_tmp176 (.Y(N1615),.A(N1464),.B(ttmp175));
OR2X1 OR_tmp177 (.Y(ttmp177),.A(N1468),.B(N1097));
OR2X1 OR_tmp178 (.Y(ttmp178),.A(N1466),.B(ttmp177));
OR2X1 OR_tmp179 (.Y(N1619),.A(N1467),.B(ttmp178));
OR2X1 OR_tmp180 (.Y(ttmp180),.A(N1471),.B(N1098));
OR2X1 OR_tmp181 (.Y(ttmp181),.A(N1469),.B(ttmp180));
OR2X1 OR_tmp182 (.Y(N1624),.A(N1470),.B(ttmp181));
OR2X1 OR_tmp183 (.Y(ttmp183),.A(N1474),.B(N1099));
OR2X1 OR_tmp184 (.Y(ttmp184),.A(N1472),.B(ttmp183));
OR2X1 OR_tmp185 (.Y(N1628),.A(N1473),.B(ttmp184));
OR2X1 OR_tmp186 (.Y(ttmp186),.A(N1477),.B(N1100));
OR2X1 OR_tmp187 (.Y(ttmp187),.A(N1475),.B(ttmp186));
OR2X1 OR_tmp188 (.Y(N1631),.A(N1476),.B(ttmp187));
OR2X1 OR_tmp189 (.Y(ttmp189),.A(N1480),.B(N1101));
OR2X1 OR_tmp190 (.Y(ttmp190),.A(N1478),.B(ttmp189));
OR2X1 OR_tmp191 (.Y(N1634),.A(N1479),.B(ttmp190));
OR2X1 OR_tmp192 (.Y(ttmp192),.A(N1483),.B(N1124));
OR2X1 OR_tmp193 (.Y(ttmp193),.A(N1481),.B(ttmp192));
OR2X1 OR_tmp194 (.Y(N1637),.A(N1482),.B(ttmp193));
OR2X1 OR_tmp195 (.Y(ttmp195),.A(N1486),.B(N1125));
OR2X1 OR_tmp196 (.Y(ttmp196),.A(N1484),.B(ttmp195));
OR2X1 OR_tmp197 (.Y(N1642),.A(N1485),.B(ttmp196));
OR2X1 OR_tmp198 (.Y(ttmp198),.A(N1489),.B(N1126));
OR2X1 OR_tmp199 (.Y(ttmp199),.A(N1487),.B(ttmp198));
OR2X1 OR_tmp200 (.Y(N1647),.A(N1488),.B(ttmp199));
OR2X1 OR_tmp201 (.Y(ttmp201),.A(N1492),.B(N1127));
OR2X1 OR_tmp202 (.Y(ttmp202),.A(N1490),.B(ttmp201));
OR2X1 OR_tmp203 (.Y(N1651),.A(N1491),.B(ttmp202));
OR2X1 OR_tmp204 (.Y(ttmp204),.A(N1495),.B(N1128));
OR2X1 OR_tmp205 (.Y(ttmp205),.A(N1493),.B(ttmp204));
OR2X1 OR_tmp206 (.Y(N1656),.A(N1494),.B(ttmp205));
OR2X1 OR_tmp207 (.Y(ttmp207),.A(N1534),.B(N1169));
OR2X1 OR_tmp208 (.Y(ttmp208),.A(N1532),.B(ttmp207));
OR2X1 OR_tmp209 (.Y(N1676),.A(N1533),.B(ttmp208));
OR2X1 OR_tmp210 (.Y(ttmp210),.A(N1537),.B(N1170));
OR2X1 OR_tmp211 (.Y(ttmp211),.A(N1535),.B(ttmp210));
OR2X1 OR_tmp212 (.Y(N1681),.A(N1536),.B(ttmp211));
OR2X1 OR_tmp213 (.Y(ttmp213),.A(N1540),.B(N1171));
OR2X1 OR_tmp214 (.Y(ttmp214),.A(N1538),.B(ttmp213));
OR2X1 OR_tmp215 (.Y(N1686),.A(N1539),.B(ttmp214));
OR2X1 OR_tmp216 (.Y(ttmp216),.A(N1543),.B(N1172));
OR2X1 OR_tmp217 (.Y(ttmp217),.A(N1541),.B(ttmp216));
OR2X1 OR_tmp218 (.Y(N1690),.A(N1542),.B(ttmp217));
OR2X1 OR_tmp219 (.Y(ttmp219),.A(N1531),.B(N1168));
OR2X1 OR_tmp220 (.Y(ttmp220),.A(N1529),.B(ttmp219));
OR2X1 OR_tmp221 (.Y(N1708),.A(N1530),.B(ttmp220));
BUFX1 BUFF1_343 (.Y(N1726),.A(N1591));
INVX1 NOT1_344 (.Y(N1770),.A(N1502));
INVX1 NOT1_345 (.Y(N1773),.A(N1506));
INVX1 NOT1_346 (.Y(N1776),.A(N1513));
INVX1 NOT1_347 (.Y(N1777),.A(N1516));
BUFX1 BUFF1_348 (.Y(N1778),.A(N1510));
BUFX1 BUFF1_349 (.Y(N1781),.A(N1510));
AND2X1 AND_tmp222 (.Y(ttmp222),.A(N1129),.B(N1513));
AND2X1 AND_tmp223 (.Y(N1784),.A(N1133),.B(ttmp222));
AND2X1 AND_tmp224 (.Y(ttmp224),.A(N1496),.B(N1516));
AND2X1 AND_tmp225 (.Y(N1785),.A(N1499),.B(ttmp224));
INVX1 NOT1_352 (.Y(N1795),.A(N1553));
INVX1 NOT1_353 (.Y(N1798),.A(N1557));
BUFX1 BUFF1_354 (.Y(N1801),.A(N1561));
BUFX1 BUFF1_355 (.Y(N1804),.A(N1561));
INVX1 NOT1_356 (.Y(N1807),.A(N1588));
INVX1 NOT1_357 (.Y(N1808),.A(N1578));
NAND2X1 NAND2_358 (.Y(N1809),.A(N1578),.B(N1581));
INVX1 NOT1_359 (.Y(N1810),.A(N1582));
INVX1 NOT1_360 (.Y(N1811),.A(N1585));
AND2X1 AND2_361 (.Y(N1813),.A(N1596),.B(N241));
AND2X1 AND2_362 (.Y(N1814),.A(N1606),.B(N241));
AND2X1 AND2_363 (.Y(N1815),.A(N1600),.B(N241));
INVX1 NOT1_364 (.Y(N1816),.A(N1642));
INVX1 NOT1_365 (.Y(N1817),.A(N1647));
INVX1 NOT1_366 (.Y(N1818),.A(N1637));
INVX1 NOT1_367 (.Y(N1819),.A(N1624));
INVX1 NOT1_368 (.Y(N1820),.A(N1619));
INVX1 NOT1_369 (.Y(N1821),.A(N1615));
AND2X1 AND_tmp226 (.Y(ttmp226),.A(N36),.B(N1591));
AND2X1 AND_tmp227 (.Y(ttmp227),.A(N496),.B(ttmp226));
AND2X1 AND_tmp228 (.Y(N1822),.A(N224),.B(ttmp227));
AND2X1 AND_tmp229 (.Y(ttmp229),.A(N1591),.B(N486));
AND2X1 AND_tmp230 (.Y(ttmp230),.A(N496),.B(ttmp229));
AND2X1 AND_tmp231 (.Y(N1823),.A(N224),.B(ttmp230));
BUFX1 BUFF1_372 (.Y(N1824),.A(N1596));
INVX1 NOT1_373 (.Y(N1827),.A(N1606));
AND2X1 AND2_374 (.Y(N1830),.A(N1600),.B(N537));
AND2X1 AND2_375 (.Y(N1831),.A(N1606),.B(N537));
AND2X1 AND2_376 (.Y(N1832),.A(N1619),.B(N246));
INVX1 NOT1_377 (.Y(N1833),.A(N1596));
INVX1 NOT1_378 (.Y(N1836),.A(N1600));
INVX1 NOT1_379 (.Y(N1841),.A(N1606));
BUFX1 BUFF1_380 (.Y(N1848),.A(N1612));
BUFX1 BUFF1_381 (.Y(N1852),.A(N1615));
BUFX1 BUFF1_382 (.Y(N1856),.A(N1619));
BUFX1 BUFF1_383 (.Y(N1863),.A(N1624));
BUFX1 BUFF1_384 (.Y(N1870),.A(N1628));
BUFX1 BUFF1_385 (.Y(N1875),.A(N1631));
BUFX1 BUFF1_386 (.Y(N1880),.A(N1634));
NAND2X1 NAND2_387 (.Y(N1885),.A(N727),.B(N1651));
NAND2X1 NAND2_388 (.Y(N1888),.A(N730),.B(N1656));
BUFX1 BUFF1_389 (.Y(N1891),.A(N1686));
AND2X1 AND2_390 (.Y(N1894),.A(N1637),.B(N425));
INVX1 NOT1_391 (.Y(N1897),.A(N1642));
AND2X1 AND_tmp232 (.Y(ttmp232),.A(N1133),.B(N1776));
AND2X1 AND_tmp233 (.Y(N1908),.A(N1496),.B(ttmp232));
AND2X1 AND_tmp234 (.Y(ttmp234),.A(N1499),.B(N1777));
AND2X1 AND_tmp235 (.Y(N1909),.A(N1129),.B(ttmp234));
AND2X1 AND2_394 (.Y(N1910),.A(N1600),.B(N637));
AND2X1 AND2_395 (.Y(N1911),.A(N1606),.B(N637));
AND2X1 AND2_396 (.Y(N1912),.A(N1612),.B(N637));
AND2X1 AND2_397 (.Y(N1913),.A(N1615),.B(N637));
AND2X1 AND2_398 (.Y(N1914),.A(N1619),.B(N643));
AND2X1 AND2_399 (.Y(N1915),.A(N1624),.B(N643));
AND2X1 AND2_400 (.Y(N1916),.A(N1628),.B(N643));
AND2X1 AND2_401 (.Y(N1917),.A(N1631),.B(N643));
AND2X1 AND2_402 (.Y(N1918),.A(N1634),.B(N643));
INVX1 NOT1_403 (.Y(N1919),.A(N1708));
AND2X1 AND2_404 (.Y(N1928),.A(N1676),.B(N693));
AND2X1 AND2_405 (.Y(N1929),.A(N1681),.B(N693));
AND2X1 AND2_406 (.Y(N1930),.A(N1686),.B(N693));
AND2X1 AND2_407 (.Y(N1931),.A(N1690),.B(N693));
AND2X1 AND2_408 (.Y(N1932),.A(N1637),.B(N699));
AND2X1 AND2_409 (.Y(N1933),.A(N1642),.B(N699));
AND2X1 AND2_410 (.Y(N1934),.A(N1647),.B(N699));
AND2X1 AND2_411 (.Y(N1935),.A(N1651),.B(N699));
BUFX1 BUFF1_412 (.Y(N1936),.A(N1600));
NAND2X1 NAND2_413 (.Y(N1939),.A(N1216),.B(N1808));
NAND2X1 NAND2_414 (.Y(N1940),.A(N1585),.B(N1810));
NAND2X1 NAND2_415 (.Y(N1941),.A(N1582),.B(N1811));
BUFX1 BUFF1_416 (.Y(N1942),.A(N1676));
BUFX1 BUFF1_417 (.Y(N1945),.A(N1686));
BUFX1 BUFF1_418 (.Y(N1948),.A(N1681));
BUFX1 BUFF1_419 (.Y(N1951),.A(N1637));
BUFX1 BUFF1_420 (.Y(N1954),.A(N1690));
BUFX1 BUFF1_421 (.Y(N1957),.A(N1647));
BUFX1 BUFF1_422 (.Y(N1960),.A(N1642));
BUFX1 BUFF1_423 (.Y(N1963),.A(N1656));
BUFX1 BUFF1_424 (.Y(N1966),.A(N1651));
OR2X1 OR2_425 (.Y(N1969),.A(N533),.B(N1815));
INVX1 NOT1_426 (.Y(N1970),.A(N1822));
INVX1 NOT1_427 (.Y(N1971),.A(N1823));
BUFX1 BUFF1_428 (.Y(N2010),.A(N1848));
BUFX1 BUFF1_429 (.Y(N2012),.A(N1852));
BUFX1 BUFF1_430 (.Y(N2014),.A(N1856));
BUFX1 BUFF1_431 (.Y(N2016),.A(N1863));
BUFX1 BUFF1_432 (.Y(N2018),.A(N1870));
BUFX1 BUFF1_433 (.Y(N2020),.A(N1875));
BUFX1 BUFF1_434 (.Y(N2022),.A(N1880));
INVX1 NOT1_435 (.Y(N2028),.A(N1778));
INVX1 NOT1_436 (.Y(N2029),.A(N1781));
NOR2X1 NOR2_437 (.Y(N2030),.A(N1908),.B(N1784));
NOR2X1 NOR2_438 (.Y(N2031),.A(N1909),.B(N1785));
AND2X1 AND_tmp236 (.Y(ttmp236),.A(N1502),.B(N1778));
AND2X1 AND_tmp237 (.Y(N2032),.A(N1506),.B(ttmp236));
AND2X1 AND_tmp238 (.Y(ttmp238),.A(N1770),.B(N1781));
AND2X1 AND_tmp239 (.Y(N2033),.A(N1773),.B(ttmp238));
OR2X1 OR2_441 (.Y(N2034),.A(N1571),.B(N1935));
INVX1 NOT1_442 (.Y(N2040),.A(N1801));
INVX1 NOT1_443 (.Y(N2041),.A(N1804));
AND2X1 AND_tmp240 (.Y(ttmp240),.A(N1553),.B(N1801));
AND2X1 AND_tmp241 (.Y(N2042),.A(N1557),.B(ttmp240));
AND2X1 AND_tmp242 (.Y(ttmp242),.A(N1795),.B(N1804));
AND2X1 AND_tmp243 (.Y(N2043),.A(N1798),.B(ttmp242));
NAND2X1 NAND2_446 (.Y(N2046),.A(N1939),.B(N1809));
NAND2X1 NAND2_447 (.Y(N2049),.A(N1940),.B(N1941));
OR2X1 OR2_448 (.Y(N2052),.A(N1544),.B(N1910));
OR2X1 OR2_449 (.Y(N2055),.A(N1545),.B(N1911));
OR2X1 OR2_450 (.Y(N2058),.A(N1546),.B(N1912));
OR2X1 OR2_451 (.Y(N2061),.A(N1547),.B(N1913));
OR2X1 OR2_452 (.Y(N2064),.A(N1548),.B(N1914));
OR2X1 OR2_453 (.Y(N2067),.A(N1549),.B(N1915));
OR2X1 OR2_454 (.Y(N2070),.A(N1550),.B(N1916));
OR2X1 OR2_455 (.Y(N2073),.A(N1551),.B(N1917));
OR2X1 OR2_456 (.Y(N2076),.A(N1552),.B(N1918));
OR2X1 OR2_457 (.Y(N2079),.A(N1564),.B(N1928));
OR2X1 OR2_458 (.Y(N2095),.A(N1565),.B(N1929));
OR2X1 OR2_459 (.Y(N2098),.A(N1566),.B(N1930));
OR2X1 OR2_460 (.Y(N2101),.A(N1567),.B(N1931));
OR2X1 OR2_461 (.Y(N2104),.A(N1568),.B(N1932));
OR2X1 OR2_462 (.Y(N2107),.A(N1569),.B(N1933));
OR2X1 OR2_463 (.Y(N2110),.A(N1570),.B(N1934));
AND2X1 AND_tmp244 (.Y(ttmp244),.A(N1894),.B(N40));
AND2X1 AND_tmp245 (.Y(N2113),.A(N1897),.B(ttmp244));
INVX1 NOT1_465 (.Y(N2119),.A(N1894));
NAND2X1 NAND2_466 (.Y(N2120),.A(N408),.B(N1827));
AND2X1 AND2_467 (.Y(N2125),.A(N1824),.B(N537));
AND2X1 AND2_468 (.Y(N2126),.A(N1852),.B(N246));
AND2X1 AND2_469 (.Y(N2127),.A(N1848),.B(N537));
INVX1 NOT1_470 (.Y(N2128),.A(N1848));
INVX1 NOT1_471 (.Y(N2135),.A(N1852));
INVX1 NOT1_472 (.Y(N2141),.A(N1863));
INVX1 NOT1_473 (.Y(N2144),.A(N1870));
INVX1 NOT1_474 (.Y(N2147),.A(N1875));
INVX1 NOT1_475 (.Y(N2150),.A(N1880));
AND2X1 AND2_476 (.Y(N2153),.A(N727),.B(N1885));
AND2X1 AND2_477 (.Y(N2154),.A(N1885),.B(N1651));
AND2X1 AND2_478 (.Y(N2155),.A(N730),.B(N1888));
AND2X1 AND2_479 (.Y(N2156),.A(N1888),.B(N1656));
AND2X1 AND_tmp246 (.Y(ttmp246),.A(N1506),.B(N2028));
AND2X1 AND_tmp247 (.Y(N2157),.A(N1770),.B(ttmp246));
AND2X1 AND_tmp248 (.Y(ttmp248),.A(N1773),.B(N2029));
AND2X1 AND_tmp249 (.Y(N2158),.A(N1502),.B(ttmp248));
INVX1 NOT1_482 (.Y(N2171),.A(N1942));
NAND2X1 NAND2_483 (.Y(N2172),.A(N1942),.B(N1919));
INVX1 NOT1_484 (.Y(N2173),.A(N1945));
INVX1 NOT1_485 (.Y(N2174),.A(N1948));
INVX1 NOT1_486 (.Y(N2175),.A(N1951));
INVX1 NOT1_487 (.Y(N2176),.A(N1954));
AND2X1 AND_tmp250 (.Y(ttmp250),.A(N1557),.B(N2040));
AND2X1 AND_tmp251 (.Y(N2177),.A(N1795),.B(ttmp250));
AND2X1 AND_tmp252 (.Y(ttmp252),.A(N1798),.B(N2041));
AND2X1 AND_tmp253 (.Y(N2178),.A(N1553),.B(ttmp252));
BUFX1 BUFF1_490 (.Y(N2185),.A(N1836));
BUFX1 BUFF1_491 (.Y(N2188),.A(N1833));
BUFX1 BUFF1_492 (.Y(N2191),.A(N1841));
INVX1 NOT1_493 (.Y(N2194),.A(N1856));
INVX1 NOT1_494 (.Y(N2197),.A(N1827));
INVX1 NOT1_495 (.Y(N2200),.A(N1936));
BUFX1 BUFF1_496 (.Y(N2201),.A(N1836));
BUFX1 BUFF1_497 (.Y(N2204),.A(N1833));
BUFX1 BUFF1_498 (.Y(N2207),.A(N1841));
BUFX1 BUFF1_499 (.Y(N2210),.A(N1824));
BUFX1 BUFF1_500 (.Y(N2213),.A(N1841));
BUFX1 BUFF1_501 (.Y(N2216),.A(N1841));
NAND2X1 NAND2_502 (.Y(N2219),.A(N2031),.B(N2030));
INVX1 NOT1_503 (.Y(N2234),.A(N1957));
INVX1 NOT1_504 (.Y(N2235),.A(N1960));
INVX1 NOT1_505 (.Y(N2236),.A(N1963));
INVX1 NOT1_506 (.Y(N2237),.A(N1966));
AND2X1 AND_tmp254 (.Y(ttmp254),.A(N1897),.B(N2119));
AND2X1 AND_tmp255 (.Y(N2250),.A(N40),.B(ttmp254));
OR2X1 OR2_508 (.Y(N2266),.A(N1831),.B(N2126));
OR2X1 OR2_509 (.Y(N2269),.A(N2127),.B(N1832));
OR2X1 OR2_510 (.Y(N2291),.A(N2153),.B(N2154));
OR2X1 OR2_511 (.Y(N2294),.A(N2155),.B(N2156));
NOR2X1 NOR2_512 (.Y(N2297),.A(N2157),.B(N2032));
NOR2X1 NOR2_513 (.Y(N2298),.A(N2158),.B(N2033));
INVX1 NOT1_514 (.Y(N2300),.A(N2046));
INVX1 NOT1_515 (.Y(N2301),.A(N2049));
NAND2X1 NAND2_516 (.Y(N2302),.A(N2052),.B(N1519));
INVX1 NOT1_517 (.Y(N2303),.A(N2052));
NAND2X1 NAND2_518 (.Y(N2304),.A(N2055),.B(N1520));
INVX1 NOT1_519 (.Y(N2305),.A(N2055));
NAND2X1 NAND2_520 (.Y(N2306),.A(N2058),.B(N1521));
INVX1 NOT1_521 (.Y(N2307),.A(N2058));
NAND2X1 NAND2_522 (.Y(N2308),.A(N2061),.B(N1522));
INVX1 NOT1_523 (.Y(N2309),.A(N2061));
NAND2X1 NAND2_524 (.Y(N2310),.A(N2064),.B(N1523));
INVX1 NOT1_525 (.Y(N2311),.A(N2064));
NAND2X1 NAND2_526 (.Y(N2312),.A(N2067),.B(N1524));
INVX1 NOT1_527 (.Y(N2313),.A(N2067));
NAND2X1 NAND2_528 (.Y(N2314),.A(N2070),.B(N1525));
INVX1 NOT1_529 (.Y(N2315),.A(N2070));
NAND2X1 NAND2_530 (.Y(N2316),.A(N2073),.B(N1526));
INVX1 NOT1_531 (.Y(N2317),.A(N2073));
NAND2X1 NAND2_532 (.Y(N2318),.A(N2076),.B(N1527));
INVX1 NOT1_533 (.Y(N2319),.A(N2076));
NAND2X1 NAND2_534 (.Y(N2320),.A(N2079),.B(N1528));
INVX1 NOT1_535 (.Y(N2321),.A(N2079));
NAND2X1 NAND2_536 (.Y(N2322),.A(N1708),.B(N2171));
NAND2X1 NAND2_537 (.Y(N2323),.A(N1948),.B(N2173));
NAND2X1 NAND2_538 (.Y(N2324),.A(N1945),.B(N2174));
NAND2X1 NAND2_539 (.Y(N2325),.A(N1954),.B(N2175));
NAND2X1 NAND2_540 (.Y(N2326),.A(N1951),.B(N2176));
NOR2X1 NOR2_541 (.Y(N2327),.A(N2177),.B(N2042));
NOR2X1 NOR2_542 (.Y(N2328),.A(N2178),.B(N2043));
NAND2X1 NAND2_543 (.Y(N2329),.A(N2095),.B(N1572));
INVX1 NOT1_544 (.Y(N2330),.A(N2095));
NAND2X1 NAND2_545 (.Y(N2331),.A(N2098),.B(N1573));
INVX1 NOT1_546 (.Y(N2332),.A(N2098));
NAND2X1 NAND2_547 (.Y(N2333),.A(N2101),.B(N1574));
INVX1 NOT1_548 (.Y(N2334),.A(N2101));
NAND2X1 NAND2_549 (.Y(N2335),.A(N2104),.B(N1575));
INVX1 NOT1_550 (.Y(N2336),.A(N2104));
NAND2X1 NAND2_551 (.Y(N2337),.A(N2107),.B(N1576));
INVX1 NOT1_552 (.Y(N2338),.A(N2107));
NAND2X1 NAND2_553 (.Y(N2339),.A(N2110),.B(N1577));
INVX1 NOT1_554 (.Y(N2340),.A(N2110));
NAND2X1 NAND2_555 (.Y(N2354),.A(N1960),.B(N2234));
NAND2X1 NAND2_556 (.Y(N2355),.A(N1957),.B(N2235));
NAND2X1 NAND2_557 (.Y(N2356),.A(N1966),.B(N2236));
NAND2X1 NAND2_558 (.Y(N2357),.A(N1963),.B(N2237));
AND2X1 AND2_559 (.Y(N2358),.A(N2120),.B(N533));
INVX1 NOT1_560 (.Y(N2359),.A(N2113));
INVX1 NOT1_561 (.Y(N2364),.A(N2185));
INVX1 NOT1_562 (.Y(N2365),.A(N2188));
INVX1 NOT1_563 (.Y(N2366),.A(N2191));
INVX1 NOT1_564 (.Y(N2367),.A(N2194));
BUFX1 BUFF1_565 (.Y(N2368),.A(N2120));
INVX1 NOT1_566 (.Y(N2372),.A(N2201));
INVX1 NOT1_567 (.Y(N2373),.A(N2204));
INVX1 NOT1_568 (.Y(N2374),.A(N2207));
INVX1 NOT1_569 (.Y(N2375),.A(N2210));
INVX1 NOT1_570 (.Y(N2376),.A(N2213));
INVX1 NOT1_571 (.Y(N2377),.A(N2113));
BUFX1 BUFF1_572 (.Y(N2382),.A(N2113));
AND2X1 AND2_573 (.Y(N2386),.A(N2120),.B(N246));
BUFX1 BUFF1_574 (.Y(N2387),.A(N2266));
BUFX1 BUFF1_575 (.Y(N2388),.A(N2266));
BUFX1 BUFF1_576 (.Y(N2389),.A(N2269));
BUFX1 BUFF1_577 (.Y(N2390),.A(N2269));
BUFX1 BUFF1_578 (.Y(N2391),.A(N2113));
INVX1 NOT1_579 (.Y(N2395),.A(N2113));
NAND2X1 NAND2_580 (.Y(N2400),.A(N2219),.B(N2300));
INVX1 NOT1_581 (.Y(N2403),.A(N2216));
INVX1 NOT1_582 (.Y(N2406),.A(N2219));
NAND2X1 NAND2_583 (.Y(N2407),.A(N1219),.B(N2303));
NAND2X1 NAND2_584 (.Y(N2408),.A(N1222),.B(N2305));
NAND2X1 NAND2_585 (.Y(N2409),.A(N1225),.B(N2307));
NAND2X1 NAND2_586 (.Y(N2410),.A(N1228),.B(N2309));
NAND2X1 NAND2_587 (.Y(N2411),.A(N1231),.B(N2311));
NAND2X1 NAND2_588 (.Y(N2412),.A(N1234),.B(N2313));
NAND2X1 NAND2_589 (.Y(N2413),.A(N1237),.B(N2315));
NAND2X1 NAND2_590 (.Y(N2414),.A(N1240),.B(N2317));
NAND2X1 NAND2_591 (.Y(N2415),.A(N1243),.B(N2319));
NAND2X1 NAND2_592 (.Y(N2416),.A(N1246),.B(N2321));
NAND2X1 NAND2_593 (.Y(N2417),.A(N2322),.B(N2172));
NAND2X1 NAND2_594 (.Y(N2421),.A(N2323),.B(N2324));
NAND2X1 NAND2_595 (.Y(N2425),.A(N2325),.B(N2326));
NAND2X1 NAND2_596 (.Y(N2428),.A(N1251),.B(N2330));
NAND2X1 NAND2_597 (.Y(N2429),.A(N1254),.B(N2332));
NAND2X1 NAND2_598 (.Y(N2430),.A(N1257),.B(N2334));
NAND2X1 NAND2_599 (.Y(N2431),.A(N1260),.B(N2336));
NAND2X1 NAND2_600 (.Y(N2432),.A(N1263),.B(N2338));
NAND2X1 NAND2_601 (.Y(N2433),.A(N1266),.B(N2340));
BUFX1 BUFF1_602 (.Y(N2434),.A(N2128));
BUFX1 BUFF1_603 (.Y(N2437),.A(N2135));
BUFX1 BUFF1_604 (.Y(N2440),.A(N2144));
BUFX1 BUFF1_605 (.Y(N2443),.A(N2141));
BUFX1 BUFF1_606 (.Y(N2446),.A(N2150));
BUFX1 BUFF1_607 (.Y(N2449),.A(N2147));
INVX1 NOT1_608 (.Y(N2452),.A(N2197));
NAND2X1 NAND2_609 (.Y(N2453),.A(N2197),.B(N2200));
BUFX1 BUFF1_610 (.Y(N2454),.A(N2128));
BUFX1 BUFF1_611 (.Y(N2457),.A(N2144));
BUFX1 BUFF1_612 (.Y(N2460),.A(N2141));
BUFX1 BUFF1_613 (.Y(N2463),.A(N2150));
BUFX1 BUFF1_614 (.Y(N2466),.A(N2147));
INVX1 NOT1_615 (.Y(N2469),.A(N2120));
BUFX1 BUFF1_616 (.Y(N2472),.A(N2128));
BUFX1 BUFF1_617 (.Y(N2475),.A(N2135));
BUFX1 BUFF1_618 (.Y(N2478),.A(N2128));
BUFX1 BUFF1_619 (.Y(N2481),.A(N2135));
NAND2X1 NAND2_620 (.Y(N2484),.A(N2298),.B(N2297));
NAND2X1 NAND2_621 (.Y(N2487),.A(N2356),.B(N2357));
NAND2X1 NAND2_622 (.Y(N2490),.A(N2354),.B(N2355));
NAND2X1 NAND2_623 (.Y(N2493),.A(N2328),.B(N2327));
OR2X1 OR2_624 (.Y(N2496),.A(N2358),.B(N1814));
NAND2X1 NAND2_625 (.Y(N2503),.A(N2188),.B(N2364));
NAND2X1 NAND2_626 (.Y(N2504),.A(N2185),.B(N2365));
NAND2X1 NAND2_627 (.Y(N2510),.A(N2204),.B(N2372));
NAND2X1 NAND2_628 (.Y(N2511),.A(N2201),.B(N2373));
OR2X1 OR2_629 (.Y(N2521),.A(N1830),.B(N2386));
NAND2X1 NAND2_630 (.Y(N2528),.A(N2046),.B(N2406));
INVX1 NOT1_631 (.Y(N2531),.A(N2291));
INVX1 NOT1_632 (.Y(N2534),.A(N2294));
BUFX1 BUFF1_633 (.Y(N2537),.A(N2250));
BUFX1 BUFF1_634 (.Y(N2540),.A(N2250));
NAND2X1 NAND2_635 (.Y(N2544),.A(N2302),.B(N2407));
NAND2X1 NAND2_636 (.Y(N2545),.A(N2304),.B(N2408));
NAND2X1 NAND2_637 (.Y(N2546),.A(N2306),.B(N2409));
NAND2X1 NAND2_638 (.Y(N2547),.A(N2308),.B(N2410));
NAND2X1 NAND2_639 (.Y(N2548),.A(N2310),.B(N2411));
NAND2X1 NAND2_640 (.Y(N2549),.A(N2312),.B(N2412));
NAND2X1 NAND2_641 (.Y(N2550),.A(N2314),.B(N2413));
NAND2X1 NAND2_642 (.Y(N2551),.A(N2316),.B(N2414));
NAND2X1 NAND2_643 (.Y(N2552),.A(N2318),.B(N2415));
NAND2X1 NAND2_644 (.Y(N2553),.A(N2320),.B(N2416));
NAND2X1 NAND2_645 (.Y(N2563),.A(N2329),.B(N2428));
NAND2X1 NAND2_646 (.Y(N2564),.A(N2331),.B(N2429));
NAND2X1 NAND2_647 (.Y(N2565),.A(N2333),.B(N2430));
NAND2X1 NAND2_648 (.Y(N2566),.A(N2335),.B(N2431));
NAND2X1 NAND2_649 (.Y(N2567),.A(N2337),.B(N2432));
NAND2X1 NAND2_650 (.Y(N2568),.A(N2339),.B(N2433));
NAND2X1 NAND2_651 (.Y(N2579),.A(N1936),.B(N2452));
BUFX1 BUFF1_652 (.Y(N2603),.A(N2359));
AND2X1 AND2_653 (.Y(N2607),.A(N1880),.B(N2377));
AND2X1 AND2_654 (.Y(N2608),.A(N1676),.B(N2377));
AND2X1 AND2_655 (.Y(N2609),.A(N1681),.B(N2377));
AND2X1 AND2_656 (.Y(N2610),.A(N1891),.B(N2377));
AND2X1 AND2_657 (.Y(N2611),.A(N1856),.B(N2382));
AND2X1 AND2_658 (.Y(N2612),.A(N1863),.B(N2382));
NAND2X1 NAND2_659 (.Y(N2613),.A(N2503),.B(N2504));
INVX1 NOT1_660 (.Y(N2617),.A(N2434));
NAND2X1 NAND2_661 (.Y(N2618),.A(N2434),.B(N2366));
NAND2X1 NAND2_662 (.Y(N2619),.A(N2437),.B(N2367));
INVX1 NOT1_663 (.Y(N2620),.A(N2437));
INVX1 NOT1_664 (.Y(N2621),.A(N2368));
NAND2X1 NAND2_665 (.Y(N2624),.A(N2510),.B(N2511));
INVX1 NOT1_666 (.Y(N2628),.A(N2454));
NAND2X1 NAND2_667 (.Y(N2629),.A(N2454),.B(N2374));
INVX1 NOT1_668 (.Y(N2630),.A(N2472));
AND2X1 AND2_669 (.Y(N2631),.A(N1856),.B(N2391));
AND2X1 AND2_670 (.Y(N2632),.A(N1863),.B(N2391));
AND2X1 AND2_671 (.Y(N2633),.A(N1880),.B(N2395));
AND2X1 AND2_672 (.Y(N2634),.A(N1676),.B(N2395));
AND2X1 AND2_673 (.Y(N2635),.A(N1681),.B(N2395));
AND2X1 AND2_674 (.Y(N2636),.A(N1891),.B(N2395));
INVX1 NOT1_675 (.Y(N2638),.A(N2382));
BUFX1 BUFF1_676 (.Y(N2643),.A(N2521));
BUFX1 BUFF1_677 (.Y(N2644),.A(N2521));
INVX1 NOT1_678 (.Y(N2645),.A(N2475));
INVX1 NOT1_679 (.Y(N2646),.A(N2391));
NAND2X1 NAND2_680 (.Y(N2652),.A(N2528),.B(N2400));
INVX1 NOT1_681 (.Y(N2655),.A(N2478));
INVX1 NOT1_682 (.Y(N2656),.A(N2481));
BUFX1 BUFF1_683 (.Y(N2659),.A(N2359));
INVX1 NOT1_684 (.Y(N2663),.A(N2484));
NAND2X1 NAND2_685 (.Y(N2664),.A(N2484),.B(N2301));
INVX1 NOT1_686 (.Y(N2665),.A(N2553));
INVX1 NOT1_687 (.Y(N2666),.A(N2552));
INVX1 NOT1_688 (.Y(N2667),.A(N2551));
INVX1 NOT1_689 (.Y(N2668),.A(N2550));
INVX1 NOT1_690 (.Y(N2669),.A(N2549));
INVX1 NOT1_691 (.Y(N2670),.A(N2548));
INVX1 NOT1_692 (.Y(N2671),.A(N2547));
INVX1 NOT1_693 (.Y(N2672),.A(N2546));
INVX1 NOT1_694 (.Y(N2673),.A(N2545));
INVX1 NOT1_695 (.Y(N2674),.A(N2544));
INVX1 NOT1_696 (.Y(N2675),.A(N2568));
INVX1 NOT1_697 (.Y(N2676),.A(N2567));
INVX1 NOT1_698 (.Y(N2677),.A(N2566));
INVX1 NOT1_699 (.Y(N2678),.A(N2565));
INVX1 NOT1_700 (.Y(N2679),.A(N2564));
INVX1 NOT1_701 (.Y(N2680),.A(N2563));
INVX1 NOT1_702 (.Y(N2681),.A(N2417));
INVX1 NOT1_703 (.Y(N2684),.A(N2421));
BUFX1 BUFF1_704 (.Y(N2687),.A(N2425));
BUFX1 BUFF1_705 (.Y(N2690),.A(N2425));
INVX1 NOT1_706 (.Y(N2693),.A(N2493));
NAND2X1 NAND2_707 (.Y(N2694),.A(N2493),.B(N1807));
INVX1 NOT1_708 (.Y(N2695),.A(N2440));
INVX1 NOT1_709 (.Y(N2696),.A(N2443));
INVX1 NOT1_710 (.Y(N2697),.A(N2446));
INVX1 NOT1_711 (.Y(N2698),.A(N2449));
INVX1 NOT1_712 (.Y(N2699),.A(N2457));
INVX1 NOT1_713 (.Y(N2700),.A(N2460));
INVX1 NOT1_714 (.Y(N2701),.A(N2463));
INVX1 NOT1_715 (.Y(N2702),.A(N2466));
NAND2X1 NAND2_716 (.Y(N2703),.A(N2579),.B(N2453));
INVX1 NOT1_717 (.Y(N2706),.A(N2469));
INVX1 NOT1_718 (.Y(N2707),.A(N2487));
INVX1 NOT1_719 (.Y(N2708),.A(N2490));
AND2X1 AND2_720 (.Y(N2709),.A(N2294),.B(N2534));
AND2X1 AND2_721 (.Y(N2710),.A(N2291),.B(N2531));
NAND2X1 NAND2_722 (.Y(N2719),.A(N2191),.B(N2617));
NAND2X1 NAND2_723 (.Y(N2720),.A(N2194),.B(N2620));
NAND2X1 NAND2_724 (.Y(N2726),.A(N2207),.B(N2628));
BUFX1 BUFF1_725 (.Y(N2729),.A(N2537));
BUFX1 BUFF1_726 (.Y(N2738),.A(N2537));
INVX1 NOT1_727 (.Y(N2743),.A(N2652));
NAND2X1 NAND2_728 (.Y(N2747),.A(N2049),.B(N2663));
AND2X1 AND_tmp256 (.Y(ttmp256),.A(N2668),.B(N2669));
AND2X1 AND_tmp257 (.Y(ttmp257),.A(N2665),.B(ttmp256));
AND2X1 AND_tmp258 (.Y(ttmp258),.A(N2666),.B(ttmp257));
AND2X1 AND_tmp259 (.Y(N2748),.A(N2667),.B(ttmp258));
AND2X1 AND_tmp260 (.Y(ttmp260),.A(N2673),.B(N2674));
AND2X1 AND_tmp261 (.Y(ttmp261),.A(N2670),.B(ttmp260));
AND2X1 AND_tmp262 (.Y(ttmp262),.A(N2671),.B(ttmp261));
AND2X1 AND_tmp263 (.Y(N2749),.A(N2672),.B(ttmp262));
AND2X1 AND2_731 (.Y(N2750),.A(N2034),.B(N2675));
AND2X1 AND_tmp264 (.Y(ttmp264),.A(N2679),.B(N2680));
AND2X1 AND_tmp265 (.Y(ttmp265),.A(N2676),.B(ttmp264));
AND2X1 AND_tmp266 (.Y(ttmp266),.A(N2677),.B(ttmp265));
AND2X1 AND_tmp267 (.Y(N2751),.A(N2678),.B(ttmp266));
NAND2X1 NAND2_733 (.Y(N2760),.A(N1588),.B(N2693));
BUFX1 BUFF1_734 (.Y(N2761),.A(N2540));
BUFX1 BUFF1_735 (.Y(N2766),.A(N2540));
NAND2X1 NAND2_736 (.Y(N2771),.A(N2443),.B(N2695));
NAND2X1 NAND2_737 (.Y(N2772),.A(N2440),.B(N2696));
NAND2X1 NAND2_738 (.Y(N2773),.A(N2449),.B(N2697));
NAND2X1 NAND2_739 (.Y(N2774),.A(N2446),.B(N2698));
NAND2X1 NAND2_740 (.Y(N2775),.A(N2460),.B(N2699));
NAND2X1 NAND2_741 (.Y(N2776),.A(N2457),.B(N2700));
NAND2X1 NAND2_742 (.Y(N2777),.A(N2466),.B(N2701));
NAND2X1 NAND2_743 (.Y(N2778),.A(N2463),.B(N2702));
NAND2X1 NAND2_744 (.Y(N2781),.A(N2490),.B(N2707));
NAND2X1 NAND2_745 (.Y(N2782),.A(N2487),.B(N2708));
OR2X1 OR2_746 (.Y(N2783),.A(N2709),.B(N2534));
OR2X1 OR2_747 (.Y(N2784),.A(N2710),.B(N2531));
AND2X1 AND2_748 (.Y(N2789),.A(N1856),.B(N2638));
AND2X1 AND2_749 (.Y(N2790),.A(N1863),.B(N2638));
AND2X1 AND2_750 (.Y(N2791),.A(N1870),.B(N2638));
AND2X1 AND2_751 (.Y(N2792),.A(N1875),.B(N2638));
INVX1 NOT1_752 (.Y(N2793),.A(N2613));
NAND2X1 NAND2_753 (.Y(N2796),.A(N2719),.B(N2618));
NAND2X1 NAND2_754 (.Y(N2800),.A(N2619),.B(N2720));
INVX1 NOT1_755 (.Y(N2803),.A(N2624));
NAND2X1 NAND2_756 (.Y(N2806),.A(N2726),.B(N2629));
AND2X1 AND2_757 (.Y(N2809),.A(N1856),.B(N2646));
AND2X1 AND2_758 (.Y(N2810),.A(N1863),.B(N2646));
AND2X1 AND2_759 (.Y(N2811),.A(N1870),.B(N2646));
AND2X1 AND2_760 (.Y(N2812),.A(N1875),.B(N2646));
AND2X1 AND2_761 (.Y(N2817),.A(N2743),.B(N14));
BUFX1 BUFF1_762 (.Y(N2820),.A(N2603));
NAND2X1 NAND2_763 (.Y(N2826),.A(N2747),.B(N2664));
AND2X1 AND2_764 (.Y(N2829),.A(N2748),.B(N2749));
AND2X1 AND2_765 (.Y(N2830),.A(N2750),.B(N2751));
BUFX1 BUFF1_766 (.Y(N2831),.A(N2659));
INVX1 NOT1_767 (.Y(N2837),.A(N2687));
INVX1 NOT1_768 (.Y(N2838),.A(N2690));
AND2X1 AND_tmp268 (.Y(ttmp268),.A(N2417),.B(N2687));
AND2X1 AND_tmp269 (.Y(N2839),.A(N2421),.B(ttmp268));
AND2X1 AND_tmp270 (.Y(ttmp270),.A(N2681),.B(N2690));
AND2X1 AND_tmp271 (.Y(N2840),.A(N2684),.B(ttmp270));
NAND2X1 NAND2_771 (.Y(N2841),.A(N2760),.B(N2694));
BUFX1 BUFF1_772 (.Y(N2844),.A(N2603));
BUFX1 BUFF1_773 (.Y(N2854),.A(N2603));
BUFX1 BUFF1_774 (.Y(N2859),.A(N2659));
BUFX1 BUFF1_775 (.Y(N2869),.A(N2659));
NAND2X1 NAND2_776 (.Y(N2874),.A(N2773),.B(N2774));
NAND2X1 NAND2_777 (.Y(N2877),.A(N2771),.B(N2772));
INVX1 NOT1_778 (.Y(N2880),.A(N2703));
NAND2X1 NAND2_779 (.Y(N2881),.A(N2703),.B(N2706));
NAND2X1 NAND2_780 (.Y(N2882),.A(N2777),.B(N2778));
NAND2X1 NAND2_781 (.Y(N2885),.A(N2775),.B(N2776));
NAND2X1 NAND2_782 (.Y(N2888),.A(N2781),.B(N2782));
NAND2X1 NAND2_783 (.Y(N2891),.A(N2783),.B(N2784));
AND2X1 AND2_784 (.Y(N2894),.A(N2607),.B(N2729));
AND2X1 AND2_785 (.Y(N2895),.A(N2608),.B(N2729));
AND2X1 AND2_786 (.Y(N2896),.A(N2609),.B(N2729));
AND2X1 AND2_787 (.Y(N2897),.A(N2610),.B(N2729));
OR2X1 OR2_788 (.Y(N2898),.A(N2789),.B(N2611));
OR2X1 OR2_789 (.Y(N2899),.A(N2790),.B(N2612));
AND2X1 AND2_790 (.Y(N2900),.A(N2791),.B(N1037));
AND2X1 AND2_791 (.Y(N2901),.A(N2792),.B(N1037));
OR2X1 OR2_792 (.Y(N2914),.A(N2809),.B(N2631));
OR2X1 OR2_793 (.Y(N2915),.A(N2810),.B(N2632));
AND2X1 AND2_794 (.Y(N2916),.A(N2811),.B(N1070));
AND2X1 AND2_795 (.Y(N2917),.A(N2812),.B(N1070));
AND2X1 AND2_796 (.Y(N2918),.A(N2633),.B(N2738));
AND2X1 AND2_797 (.Y(N2919),.A(N2634),.B(N2738));
AND2X1 AND2_798 (.Y(N2920),.A(N2635),.B(N2738));
AND2X1 AND2_799 (.Y(N2921),.A(N2636),.B(N2738));
BUFX1 BUFF1_800 (.Y(N2925),.A(N2817));
AND2X1 AND_tmp272 (.Y(ttmp272),.A(N2830),.B(N1302));
AND2X1 AND_tmp273 (.Y(N2931),.A(N2829),.B(ttmp272));
AND2X1 AND_tmp274 (.Y(ttmp274),.A(N2421),.B(N2837));
AND2X1 AND_tmp275 (.Y(N2938),.A(N2681),.B(ttmp274));
AND2X1 AND_tmp276 (.Y(ttmp276),.A(N2684),.B(N2838));
AND2X1 AND_tmp277 (.Y(N2939),.A(N2417),.B(ttmp276));
NAND2X1 NAND2_804 (.Y(N2963),.A(N2469),.B(N2880));
INVX1 NOT1_805 (.Y(N2970),.A(N2841));
INVX1 NOT1_806 (.Y(N2971),.A(N2826));
INVX1 NOT1_807 (.Y(N2972),.A(N2894));
INVX1 NOT1_808 (.Y(N2975),.A(N2895));
INVX1 NOT1_809 (.Y(N2978),.A(N2896));
INVX1 NOT1_810 (.Y(N2981),.A(N2897));
AND2X1 AND2_811 (.Y(N2984),.A(N2898),.B(N1037));
AND2X1 AND2_812 (.Y(N2985),.A(N2899),.B(N1037));
INVX1 NOT1_813 (.Y(N2986),.A(N2900));
INVX1 NOT1_814 (.Y(N2989),.A(N2901));
INVX1 NOT1_815 (.Y(N2992),.A(N2796));
BUFX1 BUFF1_816 (.Y(N2995),.A(N2800));
BUFX1 BUFF1_817 (.Y(N2998),.A(N2800));
BUFX1 BUFF1_818 (.Y(N3001),.A(N2806));
BUFX1 BUFF1_819 (.Y(N3004),.A(N2806));
AND2X1 AND2_820 (.Y(N3007),.A(N574),.B(N2820));
AND2X1 AND2_821 (.Y(N3008),.A(N2914),.B(N1070));
AND2X1 AND2_822 (.Y(N3009),.A(N2915),.B(N1070));
INVX1 NOT1_823 (.Y(N3010),.A(N2916));
INVX1 NOT1_824 (.Y(N3013),.A(N2917));
INVX1 NOT1_825 (.Y(N3016),.A(N2918));
INVX1 NOT1_826 (.Y(N3019),.A(N2919));
INVX1 NOT1_827 (.Y(N3022),.A(N2920));
INVX1 NOT1_828 (.Y(N3025),.A(N2921));
INVX1 NOT1_829 (.Y(N3028),.A(N2817));
AND2X1 AND2_830 (.Y(N3029),.A(N574),.B(N2831));
INVX1 NOT1_831 (.Y(N3030),.A(N2820));
AND2X1 AND2_832 (.Y(N3035),.A(N578),.B(N2820));
AND2X1 AND2_833 (.Y(N3036),.A(N655),.B(N2820));
AND2X1 AND2_834 (.Y(N3037),.A(N659),.B(N2820));
BUFX1 BUFF1_835 (.Y(N3038),.A(N2931));
INVX1 NOT1_836 (.Y(N3039),.A(N2831));
AND2X1 AND2_837 (.Y(N3044),.A(N578),.B(N2831));
AND2X1 AND2_838 (.Y(N3045),.A(N655),.B(N2831));
AND2X1 AND2_839 (.Y(N3046),.A(N659),.B(N2831));
NOR2X1 NOR2_840 (.Y(N3047),.A(N2938),.B(N2839));
NOR2X1 NOR2_841 (.Y(N3048),.A(N2939),.B(N2840));
INVX1 NOT1_842 (.Y(N3049),.A(N2888));
INVX1 NOT1_843 (.Y(N3050),.A(N2844));
AND2X1 AND2_844 (.Y(N3053),.A(N663),.B(N2844));
AND2X1 AND2_845 (.Y(N3054),.A(N667),.B(N2844));
AND2X1 AND2_846 (.Y(N3055),.A(N671),.B(N2844));
AND2X1 AND2_847 (.Y(N3056),.A(N675),.B(N2844));
AND2X1 AND2_848 (.Y(N3057),.A(N679),.B(N2854));
AND2X1 AND2_849 (.Y(N3058),.A(N683),.B(N2854));
AND2X1 AND2_850 (.Y(N3059),.A(N687),.B(N2854));
AND2X1 AND2_851 (.Y(N3060),.A(N705),.B(N2854));
INVX1 NOT1_852 (.Y(N3061),.A(N2859));
AND2X1 AND2_853 (.Y(N3064),.A(N663),.B(N2859));
AND2X1 AND2_854 (.Y(N3065),.A(N667),.B(N2859));
AND2X1 AND2_855 (.Y(N3066),.A(N671),.B(N2859));
AND2X1 AND2_856 (.Y(N3067),.A(N675),.B(N2859));
AND2X1 AND2_857 (.Y(N3068),.A(N679),.B(N2869));
AND2X1 AND2_858 (.Y(N3069),.A(N683),.B(N2869));
AND2X1 AND2_859 (.Y(N3070),.A(N687),.B(N2869));
AND2X1 AND2_860 (.Y(N3071),.A(N705),.B(N2869));
INVX1 NOT1_861 (.Y(N3072),.A(N2874));
INVX1 NOT1_862 (.Y(N3073),.A(N2877));
INVX1 NOT1_863 (.Y(N3074),.A(N2882));
INVX1 NOT1_864 (.Y(N3075),.A(N2885));
NAND2X1 NAND2_865 (.Y(N3076),.A(N2881),.B(N2963));
INVX1 NOT1_866 (.Y(N3079),.A(N2931));
INVX1 NOT1_867 (.Y(N3088),.A(N2984));
INVX1 NOT1_868 (.Y(N3091),.A(N2985));
INVX1 NOT1_869 (.Y(N3110),.A(N3008));
INVX1 NOT1_870 (.Y(N3113),.A(N3009));
AND2X1 AND2_871 (.Y(N3137),.A(N3055),.B(N1190));
AND2X1 AND2_872 (.Y(N3140),.A(N3056),.B(N1190));
AND2X1 AND2_873 (.Y(N3143),.A(N3057),.B(N2761));
AND2X1 AND2_874 (.Y(N3146),.A(N3058),.B(N2761));
AND2X1 AND2_875 (.Y(N3149),.A(N3059),.B(N2761));
AND2X1 AND2_876 (.Y(N3152),.A(N3060),.B(N2761));
AND2X1 AND2_877 (.Y(N3157),.A(N3066),.B(N1195));
AND2X1 AND2_878 (.Y(N3160),.A(N3067),.B(N1195));
AND2X1 AND2_879 (.Y(N3163),.A(N3068),.B(N2766));
AND2X1 AND2_880 (.Y(N3166),.A(N3069),.B(N2766));
AND2X1 AND2_881 (.Y(N3169),.A(N3070),.B(N2766));
AND2X1 AND2_882 (.Y(N3172),.A(N3071),.B(N2766));
NAND2X1 NAND2_883 (.Y(N3175),.A(N2877),.B(N3072));
NAND2X1 NAND2_884 (.Y(N3176),.A(N2874),.B(N3073));
NAND2X1 NAND2_885 (.Y(N3177),.A(N2885),.B(N3074));
NAND2X1 NAND2_886 (.Y(N3178),.A(N2882),.B(N3075));
NAND2X1 NAND2_887 (.Y(N3180),.A(N3048),.B(N3047));
INVX1 NOT1_888 (.Y(N3187),.A(N2995));
INVX1 NOT1_889 (.Y(N3188),.A(N2998));
INVX1 NOT1_890 (.Y(N3189),.A(N3001));
INVX1 NOT1_891 (.Y(N3190),.A(N3004));
AND2X1 AND_tmp278 (.Y(ttmp278),.A(N2613),.B(N2995));
AND2X1 AND_tmp279 (.Y(N3191),.A(N2796),.B(ttmp278));
AND2X1 AND_tmp280 (.Y(ttmp280),.A(N2793),.B(N2998));
AND2X1 AND_tmp281 (.Y(N3192),.A(N2992),.B(ttmp280));
AND2X1 AND_tmp282 (.Y(ttmp282),.A(N2368),.B(N3001));
AND2X1 AND_tmp283 (.Y(N3193),.A(N2624),.B(ttmp282));
AND2X1 AND_tmp284 (.Y(ttmp284),.A(N2621),.B(N3004));
AND2X1 AND_tmp285 (.Y(N3194),.A(N2803),.B(ttmp284));
NAND2X1 NAND2_896 (.Y(N3195),.A(N3076),.B(N2375));
INVX1 NOT1_897 (.Y(N3196),.A(N3076));
AND2X1 AND2_898 (.Y(N3197),.A(N687),.B(N3030));
AND2X1 AND2_899 (.Y(N3208),.A(N687),.B(N3039));
AND2X1 AND2_900 (.Y(N3215),.A(N705),.B(N3030));
AND2X1 AND2_901 (.Y(N3216),.A(N711),.B(N3030));
AND2X1 AND2_902 (.Y(N3217),.A(N715),.B(N3030));
AND2X1 AND2_903 (.Y(N3218),.A(N705),.B(N3039));
AND2X1 AND2_904 (.Y(N3219),.A(N711),.B(N3039));
AND2X1 AND2_905 (.Y(N3220),.A(N715),.B(N3039));
AND2X1 AND2_906 (.Y(N3222),.A(N719),.B(N3050));
AND2X1 AND2_907 (.Y(N3223),.A(N723),.B(N3050));
AND2X1 AND2_908 (.Y(N3230),.A(N719),.B(N3061));
AND2X1 AND2_909 (.Y(N3231),.A(N723),.B(N3061));
NAND2X1 NAND2_910 (.Y(N3238),.A(N3175),.B(N3176));
NAND2X1 NAND2_911 (.Y(N3241),.A(N3177),.B(N3178));
BUFX1 BUFF1_912 (.Y(N3244),.A(N2981));
BUFX1 BUFF1_913 (.Y(N3247),.A(N2978));
BUFX1 BUFF1_914 (.Y(N3250),.A(N2975));
BUFX1 BUFF1_915 (.Y(N3253),.A(N2972));
BUFX1 BUFF1_916 (.Y(N3256),.A(N2989));
BUFX1 BUFF1_917 (.Y(N3259),.A(N2986));
BUFX1 BUFF1_918 (.Y(N3262),.A(N3025));
BUFX1 BUFF1_919 (.Y(N3265),.A(N3022));
BUFX1 BUFF1_920 (.Y(N3268),.A(N3019));
BUFX1 BUFF1_921 (.Y(N3271),.A(N3016));
BUFX1 BUFF1_922 (.Y(N3274),.A(N3013));
BUFX1 BUFF1_923 (.Y(N3277),.A(N3010));
AND2X1 AND_tmp286 (.Y(ttmp286),.A(N2796),.B(N3187));
AND2X1 AND_tmp287 (.Y(N3281),.A(N2793),.B(ttmp286));
AND2X1 AND_tmp288 (.Y(ttmp288),.A(N2992),.B(N3188));
AND2X1 AND_tmp289 (.Y(N3282),.A(N2613),.B(ttmp288));
AND2X1 AND_tmp290 (.Y(ttmp290),.A(N2624),.B(N3189));
AND2X1 AND_tmp291 (.Y(N3283),.A(N2621),.B(ttmp290));
AND2X1 AND_tmp292 (.Y(ttmp292),.A(N2803),.B(N3190));
AND2X1 AND_tmp293 (.Y(N3284),.A(N2368),.B(ttmp292));
NAND2X1 NAND2_928 (.Y(N3286),.A(N2210),.B(N3196));
OR2X1 OR2_929 (.Y(N3288),.A(N3197),.B(N3007));
NAND2X1 NAND2_930 (.Y(N3289),.A(N3180),.B(N3049));
AND2X1 AND2_931 (.Y(N3291),.A(N3152),.B(N2981));
AND2X1 AND2_932 (.Y(N3293),.A(N3149),.B(N2978));
AND2X1 AND2_933 (.Y(N3295),.A(N3146),.B(N2975));
AND2X1 AND2_934 (.Y(N3296),.A(N2972),.B(N3143));
AND2X1 AND2_935 (.Y(N3299),.A(N3140),.B(N2989));
AND2X1 AND2_936 (.Y(N3301),.A(N3137),.B(N2986));
OR2X1 OR2_937 (.Y(N3302),.A(N3208),.B(N3029));
AND2X1 AND2_938 (.Y(N3304),.A(N3172),.B(N3025));
AND2X1 AND2_939 (.Y(N3306),.A(N3169),.B(N3022));
AND2X1 AND2_940 (.Y(N3308),.A(N3166),.B(N3019));
AND2X1 AND2_941 (.Y(N3309),.A(N3016),.B(N3163));
AND2X1 AND2_942 (.Y(N3312),.A(N3160),.B(N3013));
AND2X1 AND2_943 (.Y(N3314),.A(N3157),.B(N3010));
OR2X1 OR2_944 (.Y(N3315),.A(N3215),.B(N3035));
OR2X1 OR2_945 (.Y(N3318),.A(N3216),.B(N3036));
OR2X1 OR2_946 (.Y(N3321),.A(N3217),.B(N3037));
OR2X1 OR2_947 (.Y(N3324),.A(N3218),.B(N3044));
OR2X1 OR2_948 (.Y(N3327),.A(N3219),.B(N3045));
OR2X1 OR2_949 (.Y(N3330),.A(N3220),.B(N3046));
INVX1 NOT1_950 (.Y(N3333),.A(N3180));
OR2X1 OR2_951 (.Y(N3334),.A(N3222),.B(N3053));
OR2X1 OR2_952 (.Y(N3335),.A(N3223),.B(N3054));
OR2X1 OR2_953 (.Y(N3336),.A(N3230),.B(N3064));
OR2X1 OR2_954 (.Y(N3337),.A(N3231),.B(N3065));
BUFX1 BUFF1_955 (.Y(N3340),.A(N3152));
BUFX1 BUFF1_956 (.Y(N3344),.A(N3149));
BUFX1 BUFF1_957 (.Y(N3348),.A(N3146));
BUFX1 BUFF1_958 (.Y(N3352),.A(N3143));
BUFX1 BUFF1_959 (.Y(N3356),.A(N3140));
BUFX1 BUFF1_960 (.Y(N3360),.A(N3137));
BUFX1 BUFF1_961 (.Y(N3364),.A(N3091));
BUFX1 BUFF1_962 (.Y(N3367),.A(N3088));
BUFX1 BUFF1_963 (.Y(N3370),.A(N3172));
BUFX1 BUFF1_964 (.Y(N3374),.A(N3169));
BUFX1 BUFF1_965 (.Y(N3378),.A(N3166));
BUFX1 BUFF1_966 (.Y(N3382),.A(N3163));
BUFX1 BUFF1_967 (.Y(N3386),.A(N3160));
BUFX1 BUFF1_968 (.Y(N3390),.A(N3157));
BUFX1 BUFF1_969 (.Y(N3394),.A(N3113));
BUFX1 BUFF1_970 (.Y(N3397),.A(N3110));
NAND2X1 NAND2_971 (.Y(N3400),.A(N3195),.B(N3286));
NOR2X1 NOR2_972 (.Y(N3401),.A(N3281),.B(N3191));
NOR2X1 NOR2_973 (.Y(N3402),.A(N3282),.B(N3192));
NOR2X1 NOR2_974 (.Y(N3403),.A(N3283),.B(N3193));
NOR2X1 NOR2_975 (.Y(N3404),.A(N3284),.B(N3194));
INVX1 NOT1_976 (.Y(N3405),.A(N3238));
INVX1 NOT1_977 (.Y(N3406),.A(N3241));
AND2X1 AND2_978 (.Y(N3409),.A(N3288),.B(N1836));
NAND2X1 NAND2_979 (.Y(N3410),.A(N2888),.B(N3333));
INVX1 NOT1_980 (.Y(N3412),.A(N3244));
INVX1 NOT1_981 (.Y(N3414),.A(N3247));
INVX1 NOT1_982 (.Y(N3416),.A(N3250));
INVX1 NOT1_983 (.Y(N3418),.A(N3253));
INVX1 NOT1_984 (.Y(N3420),.A(N3256));
INVX1 NOT1_985 (.Y(N3422),.A(N3259));
AND2X1 AND2_986 (.Y(N3428),.A(N3302),.B(N1836));
INVX1 NOT1_987 (.Y(N3430),.A(N3262));
INVX1 NOT1_988 (.Y(N3432),.A(N3265));
INVX1 NOT1_989 (.Y(N3434),.A(N3268));
INVX1 NOT1_990 (.Y(N3436),.A(N3271));
INVX1 NOT1_991 (.Y(N3438),.A(N3274));
INVX1 NOT1_992 (.Y(N3440),.A(N3277));
AND2X1 AND2_993 (.Y(N3450),.A(N3334),.B(N1190));
AND2X1 AND2_994 (.Y(N3453),.A(N3335),.B(N1190));
AND2X1 AND2_995 (.Y(N3456),.A(N3336),.B(N1195));
AND2X1 AND2_996 (.Y(N3459),.A(N3337),.B(N1195));
AND2X1 AND2_997 (.Y(N3478),.A(N3400),.B(N533));
AND2X1 AND2_998 (.Y(N3479),.A(N3318),.B(N2128));
AND2X1 AND2_999 (.Y(N3480),.A(N3315),.B(N1841));
NAND2X1 NAND2_1000 (.Y(N3481),.A(N3410),.B(N3289));
INVX1 NOT1_1001 (.Y(N3482),.A(N3340));
NAND2X1 NAND2_1002 (.Y(N3483),.A(N3340),.B(N3412));
INVX1 NOT1_1003 (.Y(N3484),.A(N3344));
NAND2X1 NAND2_1004 (.Y(N3485),.A(N3344),.B(N3414));
INVX1 NOT1_1005 (.Y(N3486),.A(N3348));
NAND2X1 NAND2_1006 (.Y(N3487),.A(N3348),.B(N3416));
INVX1 NOT1_1007 (.Y(N3488),.A(N3352));
NAND2X1 NAND2_1008 (.Y(N3489),.A(N3352),.B(N3418));
INVX1 NOT1_1009 (.Y(N3490),.A(N3356));
NAND2X1 NAND2_1010 (.Y(N3491),.A(N3356),.B(N3420));
INVX1 NOT1_1011 (.Y(N3492),.A(N3360));
NAND2X1 NAND2_1012 (.Y(N3493),.A(N3360),.B(N3422));
INVX1 NOT1_1013 (.Y(N3494),.A(N3364));
INVX1 NOT1_1014 (.Y(N3496),.A(N3367));
AND2X1 AND2_1015 (.Y(N3498),.A(N3321),.B(N2135));
AND2X1 AND2_1016 (.Y(N3499),.A(N3327),.B(N2128));
AND2X1 AND2_1017 (.Y(N3500),.A(N3324),.B(N1841));
INVX1 NOT1_1018 (.Y(N3501),.A(N3370));
NAND2X1 NAND2_1019 (.Y(N3502),.A(N3370),.B(N3430));
INVX1 NOT1_1020 (.Y(N3503),.A(N3374));
NAND2X1 NAND2_1021 (.Y(N3504),.A(N3374),.B(N3432));
INVX1 NOT1_1022 (.Y(N3505),.A(N3378));
NAND2X1 NAND2_1023 (.Y(N3506),.A(N3378),.B(N3434));
INVX1 NOT1_1024 (.Y(N3507),.A(N3382));
NAND2X1 NAND2_1025 (.Y(N3508),.A(N3382),.B(N3436));
INVX1 NOT1_1026 (.Y(N3509),.A(N3386));
NAND2X1 NAND2_1027 (.Y(N3510),.A(N3386),.B(N3438));
INVX1 NOT1_1028 (.Y(N3511),.A(N3390));
NAND2X1 NAND2_1029 (.Y(N3512),.A(N3390),.B(N3440));
INVX1 NOT1_1030 (.Y(N3513),.A(N3394));
INVX1 NOT1_1031 (.Y(N3515),.A(N3397));
AND2X1 AND2_1032 (.Y(N3517),.A(N3330),.B(N2135));
NAND2X1 NAND2_1033 (.Y(N3522),.A(N3402),.B(N3401));
NAND2X1 NAND2_1034 (.Y(N3525),.A(N3404),.B(N3403));
BUFX1 BUFF1_1035 (.Y(N3528),.A(N3318));
BUFX1 BUFF1_1036 (.Y(N3531),.A(N3315));
BUFX1 BUFF1_1037 (.Y(N3534),.A(N3321));
BUFX1 BUFF1_1038 (.Y(N3537),.A(N3327));
BUFX1 BUFF1_1039 (.Y(N3540),.A(N3324));
BUFX1 BUFF1_1040 (.Y(N3543),.A(N3330));
OR2X1 OR2_1041 (.Y(N3546),.A(N3478),.B(N1813));
INVX1 NOT1_1042 (.Y(N3551),.A(N3481));
NAND2X1 NAND2_1043 (.Y(N3552),.A(N3244),.B(N3482));
NAND2X1 NAND2_1044 (.Y(N3553),.A(N3247),.B(N3484));
NAND2X1 NAND2_1045 (.Y(N3554),.A(N3250),.B(N3486));
NAND2X1 NAND2_1046 (.Y(N3555),.A(N3253),.B(N3488));
NAND2X1 NAND2_1047 (.Y(N3556),.A(N3256),.B(N3490));
NAND2X1 NAND2_1048 (.Y(N3557),.A(N3259),.B(N3492));
AND2X1 AND2_1049 (.Y(N3558),.A(N3453),.B(N3091));
AND2X1 AND2_1050 (.Y(N3559),.A(N3450),.B(N3088));
NAND2X1 NAND2_1051 (.Y(N3563),.A(N3262),.B(N3501));
NAND2X1 NAND2_1052 (.Y(N3564),.A(N3265),.B(N3503));
NAND2X1 NAND2_1053 (.Y(N3565),.A(N3268),.B(N3505));
NAND2X1 NAND2_1054 (.Y(N3566),.A(N3271),.B(N3507));
NAND2X1 NAND2_1055 (.Y(N3567),.A(N3274),.B(N3509));
NAND2X1 NAND2_1056 (.Y(N3568),.A(N3277),.B(N3511));
AND2X1 AND2_1057 (.Y(N3569),.A(N3459),.B(N3113));
AND2X1 AND2_1058 (.Y(N3570),.A(N3456),.B(N3110));
BUFX1 BUFF1_1059 (.Y(N3576),.A(N3453));
BUFX1 BUFF1_1060 (.Y(N3579),.A(N3450));
BUFX1 BUFF1_1061 (.Y(N3585),.A(N3459));
BUFX1 BUFF1_1062 (.Y(N3588),.A(N3456));
INVX1 NOT1_1063 (.Y(N3592),.A(N3522));
NAND2X1 NAND2_1064 (.Y(N3593),.A(N3522),.B(N3405));
INVX1 NOT1_1065 (.Y(N3594),.A(N3525));
NAND2X1 NAND2_1066 (.Y(N3595),.A(N3525),.B(N3406));
INVX1 NOT1_1067 (.Y(N3596),.A(N3528));
NAND2X1 NAND2_1068 (.Y(N3597),.A(N3528),.B(N2630));
NAND2X1 NAND2_1069 (.Y(N3598),.A(N3531),.B(N2376));
INVX1 NOT1_1070 (.Y(N3599),.A(N3531));
AND2X1 AND2_1071 (.Y(N3600),.A(N3551),.B(N800));
NAND2X1 NAND2_1072 (.Y(N3603),.A(N3552),.B(N3483));
NAND2X1 NAND2_1073 (.Y(N3608),.A(N3553),.B(N3485));
NAND2X1 NAND2_1074 (.Y(N3612),.A(N3554),.B(N3487));
NAND2X1 NAND2_1075 (.Y(N3615),.A(N3555),.B(N3489));
NAND2X1 NAND2_1076 (.Y(N3616),.A(N3556),.B(N3491));
NAND2X1 NAND2_1077 (.Y(N3622),.A(N3557),.B(N3493));
INVX1 NOT1_1078 (.Y(N3629),.A(N3534));
NAND2X1 NAND2_1079 (.Y(N3630),.A(N3534),.B(N2645));
INVX1 NOT1_1080 (.Y(N3631),.A(N3537));
NAND2X1 NAND2_1081 (.Y(N3632),.A(N3537),.B(N2655));
NAND2X1 NAND2_1082 (.Y(N3633),.A(N3540),.B(N2403));
INVX1 NOT1_1083 (.Y(N3634),.A(N3540));
NAND2X1 NAND2_1084 (.Y(N3635),.A(N3563),.B(N3502));
NAND2X1 NAND2_1085 (.Y(N3640),.A(N3564),.B(N3504));
NAND2X1 NAND2_1086 (.Y(N3644),.A(N3565),.B(N3506));
NAND2X1 NAND2_1087 (.Y(N3647),.A(N3566),.B(N3508));
NAND2X1 NAND2_1088 (.Y(N3648),.A(N3567),.B(N3510));
NAND2X1 NAND2_1089 (.Y(N3654),.A(N3568),.B(N3512));
INVX1 NOT1_1090 (.Y(N3661),.A(N3543));
NAND2X1 NAND2_1091 (.Y(N3662),.A(N3543),.B(N2656));
NAND2X1 NAND2_1092 (.Y(N3667),.A(N3238),.B(N3592));
NAND2X1 NAND2_1093 (.Y(N3668),.A(N3241),.B(N3594));
NAND2X1 NAND2_1094 (.Y(N3669),.A(N2472),.B(N3596));
NAND2X1 NAND2_1095 (.Y(N3670),.A(N2213),.B(N3599));
BUFX1 BUFF1_1096 (.Y(N3671),.A(N3600));
INVX1 NOT1_1097 (.Y(N3691),.A(N3576));
NAND2X1 NAND2_1098 (.Y(N3692),.A(N3576),.B(N3494));
INVX1 NOT1_1099 (.Y(N3693),.A(N3579));
NAND2X1 NAND2_1100 (.Y(N3694),.A(N3579),.B(N3496));
NAND2X1 NAND2_1101 (.Y(N3695),.A(N2475),.B(N3629));
NAND2X1 NAND2_1102 (.Y(N3696),.A(N2478),.B(N3631));
NAND2X1 NAND2_1103 (.Y(N3697),.A(N2216),.B(N3634));
INVX1 NOT1_1104 (.Y(N3716),.A(N3585));
NAND2X1 NAND2_1105 (.Y(N3717),.A(N3585),.B(N3513));
INVX1 NOT1_1106 (.Y(N3718),.A(N3588));
NAND2X1 NAND2_1107 (.Y(N3719),.A(N3588),.B(N3515));
NAND2X1 NAND2_1108 (.Y(N3720),.A(N2481),.B(N3661));
NAND2X1 NAND2_1109 (.Y(N3721),.A(N3667),.B(N3593));
NAND2X1 NAND2_1110 (.Y(N3722),.A(N3668),.B(N3595));
NAND2X1 NAND2_1111 (.Y(N3723),.A(N3669),.B(N3597));
NAND2X1 NAND2_1112 (.Y(N3726),.A(N3670),.B(N3598));
INVX1 NOT1_1113 (.Y(N3727),.A(N3600));
NAND2X1 NAND2_1114 (.Y(N3728),.A(N3364),.B(N3691));
NAND2X1 NAND2_1115 (.Y(N3729),.A(N3367),.B(N3693));
NAND2X1 NAND2_1116 (.Y(N3730),.A(N3695),.B(N3630));
AND2X1 AND_tmp294 (.Y(ttmp294),.A(N3612),.B(N3603));
AND2X1 AND_tmp295 (.Y(ttmp295),.A(N3608),.B(ttmp294));
AND2X1 AND_tmp296 (.Y(N3731),.A(N3615),.B(ttmp295));
AND2X1 AND2_1118 (.Y(N3732),.A(N3603),.B(N3293));
AND2X1 AND_tmp297 (.Y(ttmp297),.A(N3603),.B(N3295));
AND2X1 AND_tmp298 (.Y(N3733),.A(N3608),.B(ttmp297));
AND2X1 AND_tmp299 (.Y(ttmp299),.A(N3296),.B(N3608));
AND2X1 AND_tmp300 (.Y(ttmp300),.A(N3612),.B(ttmp299));
AND2X1 AND_tmp301 (.Y(N3734),.A(N3603),.B(ttmp300));
AND2X1 AND2_1121 (.Y(N3735),.A(N3616),.B(N3301));
AND2X1 AND_tmp302 (.Y(ttmp302),.A(N3616),.B(N3558));
AND2X1 AND_tmp303 (.Y(N3736),.A(N3622),.B(ttmp302));
NAND2X1 NAND2_1123 (.Y(N3737),.A(N3696),.B(N3632));
NAND2X1 NAND2_1124 (.Y(N3740),.A(N3697),.B(N3633));
NAND2X1 NAND2_1125 (.Y(N3741),.A(N3394),.B(N3716));
NAND2X1 NAND2_1126 (.Y(N3742),.A(N3397),.B(N3718));
NAND2X1 NAND2_1127 (.Y(N3743),.A(N3720),.B(N3662));
AND2X1 AND_tmp304 (.Y(ttmp304),.A(N3644),.B(N3635));
AND2X1 AND_tmp305 (.Y(ttmp305),.A(N3640),.B(ttmp304));
AND2X1 AND_tmp306 (.Y(N3744),.A(N3647),.B(ttmp305));
AND2X1 AND2_1129 (.Y(N3745),.A(N3635),.B(N3306));
AND2X1 AND_tmp307 (.Y(ttmp307),.A(N3635),.B(N3308));
AND2X1 AND_tmp308 (.Y(N3746),.A(N3640),.B(ttmp307));
AND2X1 AND_tmp309 (.Y(ttmp309),.A(N3309),.B(N3640));
AND2X1 AND_tmp310 (.Y(ttmp310),.A(N3644),.B(ttmp309));
AND2X1 AND_tmp311 (.Y(N3747),.A(N3635),.B(ttmp310));
AND2X1 AND2_1132 (.Y(N3748),.A(N3648),.B(N3314));
AND2X1 AND_tmp312 (.Y(ttmp312),.A(N3648),.B(N3569));
AND2X1 AND_tmp313 (.Y(N3749),.A(N3654),.B(ttmp312));
INVX1 NOT1_1134 (.Y(N3750),.A(N3721));
AND2X1 AND2_1135 (.Y(N3753),.A(N3722),.B(N246));
NAND2X1 NAND2_1136 (.Y(N3754),.A(N3728),.B(N3692));
NAND2X1 NAND2_1137 (.Y(N3758),.A(N3729),.B(N3694));
INVX1 NOT1_1138 (.Y(N3761),.A(N3731));
OR2X1 OR_tmp314 (.Y(ttmp314),.A(N3733),.B(N3734));
OR2X1 OR_tmp315 (.Y(ttmp315),.A(N3291),.B(ttmp314));
OR2X1 OR_tmp316 (.Y(N3762),.A(N3732),.B(ttmp315));
NAND2X1 NAND2_1140 (.Y(N3767),.A(N3741),.B(N3717));
NAND2X1 NAND2_1141 (.Y(N3771),.A(N3742),.B(N3719));
INVX1 NOT1_1142 (.Y(N3774),.A(N3744));
OR2X1 OR_tmp317 (.Y(ttmp317),.A(N3746),.B(N3747));
OR2X1 OR_tmp318 (.Y(ttmp318),.A(N3304),.B(ttmp317));
OR2X1 OR_tmp319 (.Y(N3775),.A(N3745),.B(ttmp318));
AND2X1 AND2_1144 (.Y(N3778),.A(N3723),.B(N3480));
AND2X1 AND_tmp320 (.Y(ttmp320),.A(N3723),.B(N3409));
AND2X1 AND_tmp321 (.Y(N3779),.A(N3726),.B(ttmp320));
OR2X1 OR2_1146 (.Y(N3780),.A(N2125),.B(N3753));
AND2X1 AND2_1147 (.Y(N3790),.A(N3750),.B(N800));
AND2X1 AND2_1148 (.Y(N3793),.A(N3737),.B(N3500));
AND2X1 AND_tmp322 (.Y(ttmp322),.A(N3737),.B(N3428));
AND2X1 AND_tmp323 (.Y(N3794),.A(N3740),.B(ttmp322));
OR2X1 OR_tmp324 (.Y(ttmp324),.A(N3778),.B(N3779));
OR2X1 OR_tmp325 (.Y(N3802),.A(N3479),.B(ttmp324));
BUFX1 BUFF1_1151 (.Y(N3803),.A(N3780));
BUFX1 BUFF1_1152 (.Y(N3804),.A(N3780));
INVX1 NOT1_1153 (.Y(N3805),.A(N3762));
AND2X1 AND_tmp326 (.Y(ttmp326),.A(N3616),.B(N3758));
AND2X1 AND_tmp327 (.Y(ttmp327),.A(N3622),.B(ttmp326));
AND2X1 AND_tmp328 (.Y(ttmp328),.A(N3730),.B(ttmp327));
AND2X1 AND_tmp329 (.Y(N3806),.A(N3754),.B(ttmp328));
AND2X1 AND_tmp330 (.Y(ttmp330),.A(N3559),.B(N3622));
AND2X1 AND_tmp331 (.Y(ttmp331),.A(N3754),.B(ttmp330));
AND2X1 AND_tmp332 (.Y(N3807),.A(N3616),.B(ttmp331));
AND2X1 AND_tmp333 (.Y(ttmp333),.A(N3498),.B(N3622));
AND2X1 AND_tmp334 (.Y(ttmp334),.A(N3758),.B(ttmp333));
AND2X1 AND_tmp335 (.Y(ttmp335),.A(N3754),.B(ttmp334));
AND2X1 AND_tmp336 (.Y(N3808),.A(N3616),.B(ttmp335));
BUFX1 BUFF1_1157 (.Y(N3809),.A(N3790));
OR2X1 OR_tmp337 (.Y(ttmp337),.A(N3793),.B(N3794));
OR2X1 OR_tmp338 (.Y(N3811),.A(N3499),.B(ttmp337));
INVX1 NOT1_1159 (.Y(N3812),.A(N3775));
AND2X1 AND_tmp339 (.Y(ttmp339),.A(N3648),.B(N3771));
AND2X1 AND_tmp340 (.Y(ttmp340),.A(N3654),.B(ttmp339));
AND2X1 AND_tmp341 (.Y(ttmp341),.A(N3743),.B(ttmp340));
AND2X1 AND_tmp342 (.Y(N3813),.A(N3767),.B(ttmp341));
AND2X1 AND_tmp343 (.Y(ttmp343),.A(N3570),.B(N3654));
AND2X1 AND_tmp344 (.Y(ttmp344),.A(N3767),.B(ttmp343));
AND2X1 AND_tmp345 (.Y(N3814),.A(N3648),.B(ttmp344));
AND2X1 AND_tmp346 (.Y(ttmp346),.A(N3517),.B(N3654));
AND2X1 AND_tmp347 (.Y(ttmp347),.A(N3771),.B(ttmp346));
AND2X1 AND_tmp348 (.Y(ttmp348),.A(N3767),.B(ttmp347));
AND2X1 AND_tmp349 (.Y(N3815),.A(N3648),.B(ttmp348));
OR2X1 OR_tmp350 (.Y(ttmp350),.A(N3807),.B(N3808));
OR2X1 OR_tmp351 (.Y(ttmp351),.A(N3299),.B(ttmp350));
OR2X1 OR_tmp352 (.Y(ttmp352),.A(N3735),.B(ttmp351));
OR2X1 OR_tmp353 (.Y(N3816),.A(N3736),.B(ttmp352));
AND2X1 AND2_1164 (.Y(N3817),.A(N3806),.B(N3802));
NAND2X1 NAND2_1165 (.Y(N3818),.A(N3805),.B(N3761));
INVX1 NOT1_1166 (.Y(N3819),.A(N3790));
OR2X1 OR_tmp354 (.Y(ttmp354),.A(N3814),.B(N3815));
OR2X1 OR_tmp355 (.Y(ttmp355),.A(N3312),.B(ttmp354));
OR2X1 OR_tmp356 (.Y(ttmp356),.A(N3748),.B(ttmp355));
OR2X1 OR_tmp357 (.Y(N3820),.A(N3749),.B(ttmp356));
AND2X1 AND2_1168 (.Y(N3821),.A(N3813),.B(N3811));
NAND2X1 NAND2_1169 (.Y(N3822),.A(N3812),.B(N3774));
OR2X1 OR2_1170 (.Y(N3823),.A(N3816),.B(N3817));
AND2X1 AND_tmp358 (.Y(ttmp358),.A(N3819),.B(N2841));
AND2X1 AND_tmp359 (.Y(N3826),.A(N3727),.B(ttmp358));
OR2X1 OR2_1172 (.Y(N3827),.A(N3820),.B(N3821));
INVX1 NOT1_1173 (.Y(N3834),.A(N3823));
AND2X1 AND2_1174 (.Y(N3835),.A(N3818),.B(N3823));
INVX1 NOT1_1175 (.Y(N3836),.A(N3827));
AND2X1 AND2_1176 (.Y(N3837),.A(N3822),.B(N3827));
AND2X1 AND2_1177 (.Y(N3838),.A(N3762),.B(N3834));
AND2X1 AND2_1178 (.Y(N3839),.A(N3775),.B(N3836));
OR2X1 OR2_1179 (.Y(N3840),.A(N3838),.B(N3835));
OR2X1 OR2_1180 (.Y(N3843),.A(N3839),.B(N3837));
BUFX1 BUFF1_1181 (.Y(N3851),.A(N3843));
NAND2X1 NAND2_1182 (.Y(N3852),.A(N3843),.B(N3840));
AND2X1 AND2_1183 (.Y(N3857),.A(N3843),.B(N3852));
AND2X1 AND2_1184 (.Y(N3858),.A(N3852),.B(N3840));
OR2X1 OR2_1185 (.Y(N3859),.A(N3857),.B(N3858));
INVX1 NOT1_1186 (.Y(N3864),.A(N3859));
AND2X1 AND2_1187 (.Y(N3869),.A(N3859),.B(N3864));
OR2X1 OR2_1188 (.Y(N3870),.A(N3869),.B(N3864));
INVX1 NOT1_1189 (.Y(N3875),.A(N3870));
AND2X1 AND_tmp360 (.Y(ttmp360),.A(N3028),.B(N3870));
AND2X1 AND_tmp361 (.Y(N3876),.A(N2826),.B(ttmp360));
AND2X1 AND_tmp362 (.Y(ttmp362),.A(N3876),.B(N1591));
AND2X1 AND_tmp363 (.Y(N3877),.A(N3826),.B(ttmp362));
BUFX1 BUFF1_1192 (.Y(N3881),.A(N3877));
INVX1 NOT1_1193 (.Y(N3882),.A(N3877));
BUFX1 BUFF1_1194 (.Y(N143_O),.A(N143_I));
BUFX1 BUFF1_1195 (.Y(N144_O),.A(N144_I));
BUFX1 BUFF1_1196 (.Y(N145_O),.A(N145_I));
BUFX1 BUFF1_1197 (.Y(N146_O),.A(N146_I));
BUFX1 BUFF1_1198 (.Y(N147_O),.A(N147_I));
BUFX1 BUFF1_1199 (.Y(N148_O),.A(N148_I));
BUFX1 BUFF1_1200 (.Y(N149_O),.A(N149_I));
BUFX1 BUFF1_1201 (.Y(N150_O),.A(N150_I));
BUFX1 BUFF1_1202 (.Y(N151_O),.A(N151_I));
BUFX1 BUFF1_1203 (.Y(N152_O),.A(N152_I));
BUFX1 BUFF1_1204 (.Y(N153_O),.A(N153_I));
BUFX1 BUFF1_1205 (.Y(N154_O),.A(N154_I));
BUFX1 BUFF1_1206 (.Y(N155_O),.A(N155_I));
BUFX1 BUFF1_1207 (.Y(N156_O),.A(N156_I));
BUFX1 BUFF1_1208 (.Y(N157_O),.A(N157_I));
BUFX1 BUFF1_1209 (.Y(N158_O),.A(N158_I));
BUFX1 BUFF1_1210 (.Y(N159_O),.A(N159_I));
BUFX1 BUFF1_1211 (.Y(N160_O),.A(N160_I));
BUFX1 BUFF1_1212 (.Y(N161_O),.A(N161_I));
BUFX1 BUFF1_1213 (.Y(N162_O),.A(N162_I));
BUFX1 BUFF1_1214 (.Y(N163_O),.A(N163_I));
BUFX1 BUFF1_1215 (.Y(N164_O),.A(N164_I));
BUFX1 BUFF1_1216 (.Y(N165_O),.A(N165_I));
BUFX1 BUFF1_1217 (.Y(N166_O),.A(N166_I));
BUFX1 BUFF1_1218 (.Y(N167_O),.A(N167_I));
BUFX1 BUFF1_1219 (.Y(N168_O),.A(N168_I));
BUFX1 BUFF1_1220 (.Y(N169_O),.A(N169_I));
BUFX1 BUFF1_1221 (.Y(N170_O),.A(N170_I));
BUFX1 BUFF1_1222 (.Y(N171_O),.A(N171_I));
BUFX1 BUFF1_1223 (.Y(N172_O),.A(N172_I));
BUFX1 BUFF1_1224 (.Y(N173_O),.A(N173_I));
BUFX1 BUFF1_1225 (.Y(N174_O),.A(N174_I));
BUFX1 BUFF1_1226 (.Y(N175_O),.A(N175_I));
BUFX1 BUFF1_1227 (.Y(N176_O),.A(N176_I));
BUFX1 BUFF1_1228 (.Y(N177_O),.A(N177_I));
BUFX1 BUFF1_1229 (.Y(N178_O),.A(N178_I));
BUFX1 BUFF1_1230 (.Y(N179_O),.A(N179_I));
BUFX1 BUFF1_1231 (.Y(N180_O),.A(N180_I));
BUFX1 BUFF1_1232 (.Y(N181_O),.A(N181_I));
BUFX1 BUFF1_1233 (.Y(N182_O),.A(N182_I));
BUFX1 BUFF1_1234 (.Y(N183_O),.A(N183_I));
BUFX1 BUFF1_1235 (.Y(N184_O),.A(N184_I));
BUFX1 BUFF1_1236 (.Y(N185_O),.A(N185_I));
BUFX1 BUFF1_1237 (.Y(N186_O),.A(N186_I));
BUFX1 BUFF1_1238 (.Y(N187_O),.A(N187_I));
BUFX1 BUFF1_1239 (.Y(N188_O),.A(N188_I));
BUFX1 BUFF1_1240 (.Y(N189_O),.A(N189_I));
BUFX1 BUFF1_1241 (.Y(N190_O),.A(N190_I));
BUFX1 BUFF1_1242 (.Y(N191_O),.A(N191_I));
BUFX1 BUFF1_1243 (.Y(N192_O),.A(N192_I));
BUFX1 BUFF1_1244 (.Y(N193_O),.A(N193_I));
BUFX1 BUFF1_1245 (.Y(N194_O),.A(N194_I));
BUFX1 BUFF1_1246 (.Y(N195_O),.A(N195_I));
BUFX1 BUFF1_1247 (.Y(N196_O),.A(N196_I));
BUFX1 BUFF1_1248 (.Y(N197_O),.A(N197_I));
BUFX1 BUFF1_1249 (.Y(N198_O),.A(N198_I));
BUFX1 BUFF1_1250 (.Y(N199_O),.A(N199_I));
BUFX1 BUFF1_1251 (.Y(N200_O),.A(N200_I));
BUFX1 BUFF1_1252 (.Y(N201_O),.A(N201_I));
BUFX1 BUFF1_1253 (.Y(N202_O),.A(N202_I));
BUFX1 BUFF1_1254 (.Y(N203_O),.A(N203_I));
BUFX1 BUFF1_1255 (.Y(N204_O),.A(N204_I));
BUFX1 BUFF1_1256 (.Y(N205_O),.A(N205_I));
BUFX1 BUFF1_1257 (.Y(N206_O),.A(N206_I));
BUFX1 BUFF1_1258 (.Y(N207_O),.A(N207_I));
BUFX1 BUFF1_1259 (.Y(N208_O),.A(N208_I));
BUFX1 BUFF1_1260 (.Y(N209_O),.A(N209_I));
BUFX1 BUFF1_1261 (.Y(N210_O),.A(N210_I));
BUFX1 BUFF1_1262 (.Y(N211_O),.A(N211_I));
BUFX1 BUFF1_1263 (.Y(N212_O),.A(N212_I));
BUFX1 BUFF1_1264 (.Y(N213_O),.A(N213_I));
BUFX1 BUFF1_1265 (.Y(N214_O),.A(N214_I));
BUFX1 BUFF1_1266 (.Y(N215_O),.A(N215_I));
BUFX1 BUFF1_1267 (.Y(N216_O),.A(N216_I));
BUFX1 BUFF1_1268 (.Y(N217_O),.A(N217_I));
BUFX1 BUFF1_1269 (.Y(N218_O),.A(N218_I));
endmodule 