module c3540 (N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,N5360,N5361);
input N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350;
output N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,N5360,N5361;
wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,N715,N724,N727,N736,N740,N749,N753,N763,N768,N769,N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,N825,N829,N832,N835,N836,N839,N842,N845,N848,N851,N854,N858,N861,N864,N867,N870,N874,N877,N880,N883,N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,N916,N917,N920,N923,N926,N929,N932,N935,N938,N941,N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,N1315,N1322,N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1426,N1427,N1452,N1459,N1460,N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,N1508,N1509,N1510,N1511,N1512,N1520,N1562,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,N1670,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,N1694,N1714,N1715,N1718,N1721,N1722,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,N1824,N1833,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,N1878,N1879,N1880,N1883,N1884,N1885,N1888,N1889,N1890,N1893,N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1960,N1961,N1966,N1981,N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,N2068,N2073,N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,N2178,N2179,N2180,N2181,N2183,N2184,N2185,N2188,N2191,N2194,N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,N2287,N2294,N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,N2331,N2334,N2341,N2342,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,N2435,N2436,N2437,N2438,N2439,N2440,N2443,N2444,N2445,N2448,N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,N2587,N2596,N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,N2750,N2751,N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,N2970,N2973,N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,N3138,N3141,N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,N3184,N3187,N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3410,N3413,N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,N3438,N3439,N3442,N3445,N3446,N3447,N3451,N3455,N3458,N3461,N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,N3514,N3517,N3520,N3523,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3648,N3651,N3652,N3653,N3654,N3657,N3658,N3661,N3662,N3663,N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,N3696,N3697,N3700,N3703,N3704,N3705,N3706,N3707,N3708,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3731,N3734,N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,N3789,N3800,N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,N3835,N3838,N3845,N3850,N3855,N3858,N3861,N3865,N3868,N3884,N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,N3936,N3937,N3940,N3947,N3948,N3950,N3953,N3956,N3959,N3962,N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4085,N4086,N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,N4122,N4123,N4126,N4127,N4128,N4139,N4142,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,N4186,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,N4241,N4242,N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,N4284,N4287,N4291,N4295,N4296,N4299,N4303,N4304,N4305,N4310,N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,N4359,N4362,N4365,N4368,N4371,N4376,N4377,N4387,N4390,N4393,N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,N4447,N4448,N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,N4496,N4497,N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,N4527,N4528,N4529,N4530,N4531,N4534,N4537,N4540,N4545,N4549,N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,N4602,N4603,N4608,N4613,N4616,N4619,N4623,N4628,N4629,N4630,N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,N4659,N4664,N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,N4704,N4705,N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,N4730,N4733,N4740,N4743,N4747,N4748,N4749,N4750,N4753,N4754,N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,N4822,N4823,N4826,N4829,N4830,N4831,N4838,N4844,N4847,N4850,N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,N4889,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,N4925,N4926,N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,N4952,N4953,N4954,N4957,N4964,N4965,N4968,N4969,N4970,N4973,N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,N5039,N5042,N5046,N5050,N5055,N5058,N5061,N5066,N5070,N5080,N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,N5117,N5122,N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,N5183,N5184,N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,N5212,N5215,N5217,N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,N5278,N5279,N5283,N5284,N5285,N5286,N5289,N5292,N5295,N5298,N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,N5335,N5340,N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,N5358,N5359;
BUFX1 BUFF1_1 (.Y(N655),.A(N50));
INVX1 NOT1_2 (.Y(N665),.A(N50));
BUFX1 BUFF1_3 (.Y(N670),.A(N58));
INVX1 NOT1_4 (.Y(N679),.A(N58));
BUFX1 BUFF1_5 (.Y(N683),.A(N68));
INVX1 NOT1_6 (.Y(N686),.A(N68));
BUFX1 BUFF1_7 (.Y(N690),.A(N68));
BUFX1 BUFF1_8 (.Y(N699),.A(N77));
INVX1 NOT1_9 (.Y(N702),.A(N77));
BUFX1 BUFF1_10 (.Y(N706),.A(N77));
BUFX1 BUFF1_11 (.Y(N715),.A(N87));
INVX1 NOT1_12 (.Y(N724),.A(N87));
BUFX1 BUFF1_13 (.Y(N727),.A(N97));
INVX1 NOT1_14 (.Y(N736),.A(N97));
BUFX1 BUFF1_15 (.Y(N740),.A(N107));
INVX1 NOT1_16 (.Y(N749),.A(N107));
BUFX1 BUFF1_17 (.Y(N753),.A(N116));
INVX1 NOT1_18 (.Y(N763),.A(N116));
OR2X1 OR2_19 (.Y(N768),.A(N257),.B(N264));
INVX1 NOT1_20 (.Y(N769),.A(N1));
BUFX1 BUFF1_21 (.Y(N772),.A(N1));
INVX1 NOT1_22 (.Y(N779),.A(N1));
BUFX1 BUFF1_23 (.Y(N782),.A(N13));
INVX1 NOT1_24 (.Y(N786),.A(N13));
AND2X1 AND2_25 (.Y(N793),.A(N13),.B(N20));
INVX1 NOT1_26 (.Y(N794),.A(N20));
BUFX1 BUFF1_27 (.Y(N798),.A(N20));
INVX1 NOT1_28 (.Y(N803),.A(N20));
INVX1 NOT1_29 (.Y(N820),.A(N33));
BUFX1 BUFF1_30 (.Y(N821),.A(N33));
INVX1 NOT1_31 (.Y(N825),.A(N33));
AND2X1 AND2_32 (.Y(N829),.A(N33),.B(N41));
INVX1 NOT1_33 (.Y(N832),.A(N41));
OR2X1 OR2_34 (.Y(N835),.A(N41),.B(N45));
BUFX1 BUFF1_35 (.Y(N836),.A(N45));
INVX1 NOT1_36 (.Y(N839),.A(N45));
INVX1 NOT1_37 (.Y(N842),.A(N50));
BUFX1 BUFF1_38 (.Y(N845),.A(N58));
INVX1 NOT1_39 (.Y(N848),.A(N58));
BUFX1 BUFF1_40 (.Y(N851),.A(N68));
INVX1 NOT1_41 (.Y(N854),.A(N68));
BUFX1 BUFF1_42 (.Y(N858),.A(N87));
INVX1 NOT1_43 (.Y(N861),.A(N87));
BUFX1 BUFF1_44 (.Y(N864),.A(N97));
INVX1 NOT1_45 (.Y(N867),.A(N97));
INVX1 NOT1_46 (.Y(N870),.A(N107));
BUFX1 BUFF1_47 (.Y(N874),.A(N1));
BUFX1 BUFF1_48 (.Y(N877),.A(N68));
BUFX1 BUFF1_49 (.Y(N880),.A(N107));
INVX1 NOT1_50 (.Y(N883),.A(N20));
BUFX1 BUFF1_51 (.Y(N886),.A(N190));
INVX1 NOT1_52 (.Y(N889),.A(N200));
AND2X1 AND2_53 (.Y(N890),.A(N20),.B(N200));
NAND2X1 NAND2_54 (.Y(N891),.A(N20),.B(N200));
AND2X1 AND2_55 (.Y(N892),.A(N20),.B(N179));
INVX1 NOT1_56 (.Y(N895),.A(N20));
OR2X1 OR2_57 (.Y(N896),.A(N349),.B(N33));
NAND2X1 NAND2_58 (.Y(N913),.A(N1),.B(N13));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(N20),.B(N33));
NAND2X1 NAND_tmp2 (.Y(N914),.A(N1),.B(ttmp1));
INVX1 NOT1_60 (.Y(N915),.A(N20));
INVX1 NOT1_61 (.Y(N916),.A(N33));
BUFX1 BUFF1_62 (.Y(N917),.A(N179));
INVX1 NOT1_63 (.Y(N920),.A(N213));
BUFX1 BUFF1_64 (.Y(N923),.A(N343));
BUFX1 BUFF1_65 (.Y(N926),.A(N226));
BUFX1 BUFF1_66 (.Y(N929),.A(N232));
BUFX1 BUFF1_67 (.Y(N932),.A(N238));
BUFX1 BUFF1_68 (.Y(N935),.A(N244));
BUFX1 BUFF1_69 (.Y(N938),.A(N250));
BUFX1 BUFF1_70 (.Y(N941),.A(N257));
BUFX1 BUFF1_71 (.Y(N944),.A(N264));
BUFX1 BUFF1_72 (.Y(N947),.A(N270));
BUFX1 BUFF1_73 (.Y(N950),.A(N50));
BUFX1 BUFF1_74 (.Y(N953),.A(N58));
BUFX1 BUFF1_75 (.Y(N956),.A(N58));
BUFX1 BUFF1_76 (.Y(N959),.A(N97));
BUFX1 BUFF1_77 (.Y(N962),.A(N97));
BUFX1 BUFF1_78 (.Y(N965),.A(N330));
AND2X1 AND2_79 (.Y(N1067),.A(N250),.B(N768));
OR2X1 OR2_80 (.Y(N1117),.A(N820),.B(N20));
OR2X1 OR2_81 (.Y(N1179),.A(N895),.B(N169));
INVX1 NOT1_82 (.Y(N1196),.A(N793));
OR2X1 OR2_83 (.Y(N1197),.A(N915),.B(N1));
AND2X1 AND2_84 (.Y(N1202),.A(N913),.B(N914));
OR2X1 OR2_85 (.Y(N1219),.A(N916),.B(N1));
AND2X1 AND_tmp3 (.Y(ttmp3),.A(N848),.B(N854));
AND2X1 AND_tmp4 (.Y(N1250),.A(N842),.B(ttmp3));
NAND2X1 NAND2_87 (.Y(N1251),.A(N226),.B(N655));
NAND2X1 NAND2_88 (.Y(N1252),.A(N232),.B(N670));
NAND2X1 NAND2_89 (.Y(N1253),.A(N238),.B(N690));
NAND2X1 NAND2_90 (.Y(N1254),.A(N244),.B(N706));
NAND2X1 NAND2_91 (.Y(N1255),.A(N250),.B(N715));
NAND2X1 NAND2_92 (.Y(N1256),.A(N257),.B(N727));
NAND2X1 NAND2_93 (.Y(N1257),.A(N264),.B(N740));
NAND2X1 NAND2_94 (.Y(N1258),.A(N270),.B(N753));
INVX1 NOT1_95 (.Y(N1259),.A(N926));
INVX1 NOT1_96 (.Y(N1260),.A(N929));
INVX1 NOT1_97 (.Y(N1261),.A(N932));
INVX1 NOT1_98 (.Y(N1262),.A(N935));
NAND2X1 NAND2_99 (.Y(N1263),.A(N679),.B(N686));
NAND2X1 NAND2_100 (.Y(N1264),.A(N736),.B(N749));
NAND2X1 NAND2_101 (.Y(N1267),.A(N683),.B(N699));
BUFX1 BUFF1_102 (.Y(N1268),.A(N665));
INVX1 NOT1_103 (.Y(N1271),.A(N953));
INVX1 NOT1_104 (.Y(N1272),.A(N959));
BUFX1 BUFF1_105 (.Y(N1273),.A(N839));
BUFX1 BUFF1_106 (.Y(N1276),.A(N839));
BUFX1 BUFF1_107 (.Y(N1279),.A(N782));
BUFX1 BUFF1_108 (.Y(N1298),.A(N825));
BUFX1 BUFF1_109 (.Y(N1302),.A(N832));
AND2X1 AND2_110 (.Y(N1306),.A(N779),.B(N835));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(N836),.B(N832));
AND2X1 AND_tmp6 (.Y(N1315),.A(N779),.B(ttmp5));
AND2X1 AND2_112 (.Y(N1322),.A(N769),.B(N836));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(N786),.B(N798));
AND2X1 AND_tmp8 (.Y(N1325),.A(N772),.B(ttmp7));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(N786),.B(N798));
NAND2X1 NAND_tmp10 (.Y(N1328),.A(N772),.B(ttmp9));
NAND2X1 NAND2_115 (.Y(N1331),.A(N772),.B(N786));
BUFX1 BUFF1_116 (.Y(N1334),.A(N874));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(N794),.B(N45));
NAND2X1 NAND_tmp12 (.Y(N1337),.A(N782),.B(ttmp11));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(N848),.B(N854));
NAND2X1 NAND_tmp14 (.Y(N1338),.A(N842),.B(ttmp13));
INVX1 NOT1_119 (.Y(N1339),.A(N956));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(N867),.B(N870));
AND2X1 AND_tmp16 (.Y(N1340),.A(N861),.B(ttmp15));
AND2X1 AND_tmp17 (.Y(ttmp17),.A(N867),.B(N870));
NAND2X1 NAND_tmp18 (.Y(N1343),.A(N861),.B(ttmp17));
INVX1 NOT1_122 (.Y(N1344),.A(N962));
INVX1 NOT1_123 (.Y(N1345),.A(N803));
INVX1 NOT1_124 (.Y(N1346),.A(N803));
INVX1 NOT1_125 (.Y(N1347),.A(N803));
INVX1 NOT1_126 (.Y(N1348),.A(N803));
INVX1 NOT1_127 (.Y(N1349),.A(N803));
INVX1 NOT1_128 (.Y(N1350),.A(N803));
INVX1 NOT1_129 (.Y(N1351),.A(N803));
INVX1 NOT1_130 (.Y(N1352),.A(N803));
OR2X1 OR2_131 (.Y(N1353),.A(N883),.B(N886));
NOR2X1 NOR2_132 (.Y(N1358),.A(N883),.B(N886));
BUFX1 BUFF1_133 (.Y(N1363),.A(N892));
INVX1 NOT1_134 (.Y(N1366),.A(N892));
BUFX1 BUFF1_135 (.Y(N1369),.A(N821));
BUFX1 BUFF1_136 (.Y(N1384),.A(N825));
INVX1 NOT1_137 (.Y(N1401),.A(N896));
INVX1 NOT1_138 (.Y(N1402),.A(N896));
INVX1 NOT1_139 (.Y(N1403),.A(N896));
INVX1 NOT1_140 (.Y(N1404),.A(N896));
INVX1 NOT1_141 (.Y(N1405),.A(N896));
INVX1 NOT1_142 (.Y(N1406),.A(N896));
INVX1 NOT1_143 (.Y(N1407),.A(N896));
INVX1 NOT1_144 (.Y(N1408),.A(N896));
OR2X1 OR2_145 (.Y(N1409),.A(N1),.B(N1196));
INVX1 NOT1_146 (.Y(N1426),.A(N829));
INVX1 NOT1_147 (.Y(N1427),.A(N829));
AND2X1 AND_tmp19 (.Y(ttmp19),.A(N782),.B(N794));
AND2X1 AND_tmp20 (.Y(N1452),.A(N769),.B(ttmp19));
INVX1 NOT1_149 (.Y(N1459),.A(N917));
INVX1 NOT1_150 (.Y(N1460),.A(N965));
OR2X1 OR2_151 (.Y(N1461),.A(N920),.B(N923));
NOR2X1 NOR2_152 (.Y(N1464),.A(N920),.B(N923));
INVX1 NOT1_153 (.Y(N1467),.A(N938));
INVX1 NOT1_154 (.Y(N1468),.A(N941));
INVX1 NOT1_155 (.Y(N1469),.A(N944));
INVX1 NOT1_156 (.Y(N1470),.A(N947));
BUFX1 BUFF1_157 (.Y(N1471),.A(N679));
INVX1 NOT1_158 (.Y(N1474),.A(N950));
BUFX1 BUFF1_159 (.Y(N1475),.A(N686));
BUFX1 BUFF1_160 (.Y(N1478),.A(N702));
BUFX1 BUFF1_161 (.Y(N1481),.A(N724));
BUFX1 BUFF1_162 (.Y(N1484),.A(N736));
BUFX1 BUFF1_163 (.Y(N1487),.A(N749));
BUFX1 BUFF1_164 (.Y(N1490),.A(N763));
BUFX1 BUFF1_165 (.Y(N1493),.A(N877));
BUFX1 BUFF1_166 (.Y(N1496),.A(N877));
BUFX1 BUFF1_167 (.Y(N1499),.A(N880));
BUFX1 BUFF1_168 (.Y(N1502),.A(N880));
NAND2X1 NAND2_169 (.Y(N1505),.A(N702),.B(N1250));
AND2X1 AND_tmp21 (.Y(ttmp21),.A(N1253),.B(N1254));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(N1251),.B(ttmp21));
AND2X1 AND_tmp23 (.Y(N1507),.A(N1252),.B(ttmp22));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(N1257),.B(N1258));
AND2X1 AND_tmp25 (.Y(ttmp25),.A(N1255),.B(ttmp24));
AND2X1 AND_tmp26 (.Y(N1508),.A(N1256),.B(ttmp25));
NAND2X1 NAND2_172 (.Y(N1509),.A(N929),.B(N1259));
NAND2X1 NAND2_173 (.Y(N1510),.A(N926),.B(N1260));
NAND2X1 NAND2_174 (.Y(N1511),.A(N935),.B(N1261));
NAND2X1 NAND2_175 (.Y(N1512),.A(N932),.B(N1262));
AND2X1 AND2_176 (.Y(N1520),.A(N655),.B(N1263));
AND2X1 AND2_177 (.Y(N1562),.A(N874),.B(N1337));
INVX1 NOT1_178 (.Y(N1579),.A(N1117));
AND2X1 AND2_179 (.Y(N1580),.A(N803),.B(N1117));
AND2X1 AND2_180 (.Y(N1581),.A(N1338),.B(N1345));
INVX1 NOT1_181 (.Y(N1582),.A(N1117));
AND2X1 AND2_182 (.Y(N1583),.A(N803),.B(N1117));
INVX1 NOT1_183 (.Y(N1584),.A(N1117));
AND2X1 AND2_184 (.Y(N1585),.A(N803),.B(N1117));
AND2X1 AND2_185 (.Y(N1586),.A(N854),.B(N1347));
INVX1 NOT1_186 (.Y(N1587),.A(N1117));
AND2X1 AND2_187 (.Y(N1588),.A(N803),.B(N1117));
AND2X1 AND2_188 (.Y(N1589),.A(N77),.B(N1348));
INVX1 NOT1_189 (.Y(N1590),.A(N1117));
AND2X1 AND2_190 (.Y(N1591),.A(N803),.B(N1117));
AND2X1 AND2_191 (.Y(N1592),.A(N1343),.B(N1349));
INVX1 NOT1_192 (.Y(N1593),.A(N1117));
AND2X1 AND2_193 (.Y(N1594),.A(N803),.B(N1117));
INVX1 NOT1_194 (.Y(N1595),.A(N1117));
AND2X1 AND2_195 (.Y(N1596),.A(N803),.B(N1117));
AND2X1 AND2_196 (.Y(N1597),.A(N870),.B(N1351));
INVX1 NOT1_197 (.Y(N1598),.A(N1117));
AND2X1 AND2_198 (.Y(N1599),.A(N803),.B(N1117));
AND2X1 AND2_199 (.Y(N1600),.A(N116),.B(N1352));
AND2X1 AND2_200 (.Y(N1643),.A(N222),.B(N1401));
AND2X1 AND2_201 (.Y(N1644),.A(N223),.B(N1402));
AND2X1 AND2_202 (.Y(N1645),.A(N226),.B(N1403));
AND2X1 AND2_203 (.Y(N1646),.A(N232),.B(N1404));
AND2X1 AND2_204 (.Y(N1647),.A(N238),.B(N1405));
AND2X1 AND2_205 (.Y(N1648),.A(N244),.B(N1406));
AND2X1 AND2_206 (.Y(N1649),.A(N250),.B(N1407));
AND2X1 AND2_207 (.Y(N1650),.A(N257),.B(N1408));
AND2X1 AND_tmp27 (.Y(ttmp27),.A(N13),.B(N1426));
AND2X1 AND_tmp28 (.Y(N1667),.A(N1),.B(ttmp27));
AND2X1 AND_tmp29 (.Y(ttmp29),.A(N13),.B(N1427));
AND2X1 AND_tmp30 (.Y(N1670),.A(N1),.B(ttmp29));
INVX1 NOT1_210 (.Y(N1673),.A(N1202));
INVX1 NOT1_211 (.Y(N1674),.A(N1202));
INVX1 NOT1_212 (.Y(N1675),.A(N1202));
INVX1 NOT1_213 (.Y(N1676),.A(N1202));
INVX1 NOT1_214 (.Y(N1677),.A(N1202));
INVX1 NOT1_215 (.Y(N1678),.A(N1202));
INVX1 NOT1_216 (.Y(N1679),.A(N1202));
INVX1 NOT1_217 (.Y(N1680),.A(N1202));
NAND2X1 NAND2_218 (.Y(N1691),.A(N941),.B(N1467));
NAND2X1 NAND2_219 (.Y(N1692),.A(N938),.B(N1468));
NAND2X1 NAND2_220 (.Y(N1693),.A(N947),.B(N1469));
NAND2X1 NAND2_221 (.Y(N1694),.A(N944),.B(N1470));
INVX1 NOT1_222 (.Y(N1713),.A(N1505));
AND2X1 AND2_223 (.Y(N1714),.A(N87),.B(N1264));
NAND2X1 NAND2_224 (.Y(N1715),.A(N1509),.B(N1510));
NAND2X1 NAND2_225 (.Y(N1718),.A(N1511),.B(N1512));
NAND2X1 NAND2_226 (.Y(N1721),.A(N1507),.B(N1508));
AND2X1 AND2_227 (.Y(N1722),.A(N763),.B(N1340));
NAND2X1 NAND2_228 (.Y(N1725),.A(N763),.B(N1340));
INVX1 NOT1_229 (.Y(N1726),.A(N1268));
NAND2X1 NAND2_230 (.Y(N1727),.A(N1493),.B(N1271));
INVX1 NOT1_231 (.Y(N1728),.A(N1493));
AND2X1 AND2_232 (.Y(N1729),.A(N683),.B(N1268));
NAND2X1 NAND2_233 (.Y(N1730),.A(N1499),.B(N1272));
INVX1 NOT1_234 (.Y(N1731),.A(N1499));
NAND2X1 NAND2_235 (.Y(N1735),.A(N87),.B(N1264));
INVX1 NOT1_236 (.Y(N1736),.A(N1273));
INVX1 NOT1_237 (.Y(N1737),.A(N1276));
NAND2X1 NAND2_238 (.Y(N1738),.A(N1325),.B(N821));
NAND2X1 NAND2_239 (.Y(N1747),.A(N1325),.B(N825));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(N1279),.B(N798));
NAND2X1 NAND_tmp32 (.Y(N1756),.A(N772),.B(ttmp31));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(N798),.B(N1302));
AND2X1 AND_tmp34 (.Y(ttmp34),.A(N772),.B(ttmp33));
NAND2X1 NAND_tmp35 (.Y(N1761),.A(N786),.B(ttmp34));
NAND2X1 NAND2_242 (.Y(N1764),.A(N1496),.B(N1339));
INVX1 NOT1_243 (.Y(N1765),.A(N1496));
NAND2X1 NAND2_244 (.Y(N1766),.A(N1502),.B(N1344));
INVX1 NOT1_245 (.Y(N1767),.A(N1502));
INVX1 NOT1_246 (.Y(N1768),.A(N1328));
INVX1 NOT1_247 (.Y(N1769),.A(N1334));
INVX1 NOT1_248 (.Y(N1770),.A(N1331));
AND2X1 AND2_249 (.Y(N1787),.A(N845),.B(N1579));
AND2X1 AND2_250 (.Y(N1788),.A(N150),.B(N1580));
AND2X1 AND2_251 (.Y(N1789),.A(N851),.B(N1582));
AND2X1 AND2_252 (.Y(N1790),.A(N159),.B(N1583));
AND2X1 AND2_253 (.Y(N1791),.A(N77),.B(N1584));
AND2X1 AND2_254 (.Y(N1792),.A(N50),.B(N1585));
AND2X1 AND2_255 (.Y(N1793),.A(N858),.B(N1587));
AND2X1 AND2_256 (.Y(N1794),.A(N845),.B(N1588));
AND2X1 AND2_257 (.Y(N1795),.A(N864),.B(N1590));
AND2X1 AND2_258 (.Y(N1796),.A(N851),.B(N1591));
AND2X1 AND2_259 (.Y(N1797),.A(N107),.B(N1593));
AND2X1 AND2_260 (.Y(N1798),.A(N77),.B(N1594));
AND2X1 AND2_261 (.Y(N1799),.A(N116),.B(N1595));
AND2X1 AND2_262 (.Y(N1800),.A(N858),.B(N1596));
AND2X1 AND2_263 (.Y(N1801),.A(N283),.B(N1598));
AND2X1 AND2_264 (.Y(N1802),.A(N864),.B(N1599));
AND2X1 AND2_265 (.Y(N1803),.A(N200),.B(N1363));
AND2X1 AND2_266 (.Y(N1806),.A(N889),.B(N1363));
AND2X1 AND2_267 (.Y(N1809),.A(N890),.B(N1366));
AND2X1 AND2_268 (.Y(N1812),.A(N891),.B(N1366));
NAND2X1 NAND2_269 (.Y(N1815),.A(N1298),.B(N1302));
NAND2X1 NAND2_270 (.Y(N1818),.A(N821),.B(N1302));
AND2X1 AND_tmp36 (.Y(ttmp36),.A(N1279),.B(N1179));
NAND2X1 NAND_tmp37 (.Y(N1821),.A(N772),.B(ttmp36));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(N794),.B(N1298));
NAND2X1 NAND_tmp39 (.Y(N1824),.A(N786),.B(ttmp38));
NAND2X1 NAND2_273 (.Y(N1833),.A(N786),.B(N1298));
INVX1 NOT1_274 (.Y(N1842),.A(N1369));
INVX1 NOT1_275 (.Y(N1843),.A(N1369));
INVX1 NOT1_276 (.Y(N1844),.A(N1369));
INVX1 NOT1_277 (.Y(N1845),.A(N1369));
INVX1 NOT1_278 (.Y(N1846),.A(N1369));
INVX1 NOT1_279 (.Y(N1847),.A(N1369));
INVX1 NOT1_280 (.Y(N1848),.A(N1369));
INVX1 NOT1_281 (.Y(N1849),.A(N1384));
AND2X1 AND2_282 (.Y(N1850),.A(N1384),.B(N896));
INVX1 NOT1_283 (.Y(N1851),.A(N1384));
AND2X1 AND2_284 (.Y(N1852),.A(N1384),.B(N896));
INVX1 NOT1_285 (.Y(N1853),.A(N1384));
AND2X1 AND2_286 (.Y(N1854),.A(N1384),.B(N896));
INVX1 NOT1_287 (.Y(N1855),.A(N1384));
AND2X1 AND2_288 (.Y(N1856),.A(N1384),.B(N896));
INVX1 NOT1_289 (.Y(N1857),.A(N1384));
AND2X1 AND2_290 (.Y(N1858),.A(N1384),.B(N896));
INVX1 NOT1_291 (.Y(N1859),.A(N1384));
AND2X1 AND2_292 (.Y(N1860),.A(N1384),.B(N896));
INVX1 NOT1_293 (.Y(N1861),.A(N1384));
AND2X1 AND2_294 (.Y(N1862),.A(N1384),.B(N896));
INVX1 NOT1_295 (.Y(N1863),.A(N1384));
AND2X1 AND2_296 (.Y(N1864),.A(N1384),.B(N896));
AND2X1 AND2_297 (.Y(N1869),.A(N1202),.B(N1409));
NOR2X1 NOR2_298 (.Y(N1870),.A(N50),.B(N1409));
INVX1 NOT1_299 (.Y(N1873),.A(N1306));
AND2X1 AND2_300 (.Y(N1874),.A(N1202),.B(N1409));
NOR2X1 NOR2_301 (.Y(N1875),.A(N58),.B(N1409));
INVX1 NOT1_302 (.Y(N1878),.A(N1306));
AND2X1 AND2_303 (.Y(N1879),.A(N1202),.B(N1409));
NOR2X1 NOR2_304 (.Y(N1880),.A(N68),.B(N1409));
INVX1 NOT1_305 (.Y(N1883),.A(N1306));
AND2X1 AND2_306 (.Y(N1884),.A(N1202),.B(N1409));
NOR2X1 NOR2_307 (.Y(N1885),.A(N77),.B(N1409));
INVX1 NOT1_308 (.Y(N1888),.A(N1306));
AND2X1 AND2_309 (.Y(N1889),.A(N1202),.B(N1409));
NOR2X1 NOR2_310 (.Y(N1890),.A(N87),.B(N1409));
INVX1 NOT1_311 (.Y(N1893),.A(N1322));
AND2X1 AND2_312 (.Y(N1894),.A(N1202),.B(N1409));
NOR2X1 NOR2_313 (.Y(N1895),.A(N97),.B(N1409));
INVX1 NOT1_314 (.Y(N1898),.A(N1315));
AND2X1 AND2_315 (.Y(N1899),.A(N1202),.B(N1409));
NOR2X1 NOR2_316 (.Y(N1900),.A(N107),.B(N1409));
INVX1 NOT1_317 (.Y(N1903),.A(N1315));
AND2X1 AND2_318 (.Y(N1904),.A(N1202),.B(N1409));
NOR2X1 NOR2_319 (.Y(N1905),.A(N116),.B(N1409));
INVX1 NOT1_320 (.Y(N1908),.A(N1315));
AND2X1 AND2_321 (.Y(N1909),.A(N1452),.B(N213));
NAND2X1 NAND2_322 (.Y(N1912),.A(N1452),.B(N213));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(N213),.B(N343));
AND2X1 AND_tmp41 (.Y(N1913),.A(N1452),.B(ttmp40));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(N213),.B(N343));
NAND2X1 NAND_tmp43 (.Y(N1917),.A(N1452),.B(ttmp42));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(N213),.B(N343));
AND2X1 AND_tmp45 (.Y(N1922),.A(N1452),.B(ttmp44));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(N213),.B(N343));
NAND2X1 NAND_tmp47 (.Y(N1926),.A(N1452),.B(ttmp46));
BUFX1 BUFF1_327 (.Y(N1930),.A(N1464));
NAND2X1 NAND2_328 (.Y(N1933),.A(N1691),.B(N1692));
NAND2X1 NAND2_329 (.Y(N1936),.A(N1693),.B(N1694));
INVX1 NOT1_330 (.Y(N1939),.A(N1471));
NAND2X1 NAND2_331 (.Y(N1940),.A(N1471),.B(N1474));
INVX1 NOT1_332 (.Y(N1941),.A(N1475));
INVX1 NOT1_333 (.Y(N1942),.A(N1478));
INVX1 NOT1_334 (.Y(N1943),.A(N1481));
INVX1 NOT1_335 (.Y(N1944),.A(N1484));
INVX1 NOT1_336 (.Y(N1945),.A(N1487));
INVX1 NOT1_337 (.Y(N1946),.A(N1490));
INVX1 NOT1_338 (.Y(N1947),.A(N1714));
NAND2X1 NAND2_339 (.Y(N1960),.A(N953),.B(N1728));
NAND2X1 NAND2_340 (.Y(N1961),.A(N959),.B(N1731));
AND2X1 AND2_341 (.Y(N1966),.A(N1520),.B(N1276));
NAND2X1 NAND2_342 (.Y(N1981),.A(N956),.B(N1765));
NAND2X1 NAND2_343 (.Y(N1982),.A(N962),.B(N1767));
AND2X1 AND2_344 (.Y(N1983),.A(N1067),.B(N1768));
OR2X1 OR_tmp48 (.Y(ttmp48),.A(N1787),.B(N1788));
OR2X1 OR_tmp49 (.Y(N1986),.A(N1581),.B(ttmp48));
OR2X1 OR_tmp50 (.Y(ttmp50),.A(N1791),.B(N1792));
OR2X1 OR_tmp51 (.Y(N1987),.A(N1586),.B(ttmp50));
OR2X1 OR_tmp52 (.Y(ttmp52),.A(N1793),.B(N1794));
OR2X1 OR_tmp53 (.Y(N1988),.A(N1589),.B(ttmp52));
OR2X1 OR_tmp54 (.Y(ttmp54),.A(N1795),.B(N1796));
OR2X1 OR_tmp55 (.Y(N1989),.A(N1592),.B(ttmp54));
OR2X1 OR_tmp56 (.Y(ttmp56),.A(N1799),.B(N1800));
OR2X1 OR_tmp57 (.Y(N1990),.A(N1597),.B(ttmp56));
OR2X1 OR_tmp58 (.Y(ttmp58),.A(N1801),.B(N1802));
OR2X1 OR_tmp59 (.Y(N1991),.A(N1600),.B(ttmp58));
AND2X1 AND2_351 (.Y(N2022),.A(N77),.B(N1849));
AND2X1 AND2_352 (.Y(N2023),.A(N223),.B(N1850));
AND2X1 AND2_353 (.Y(N2024),.A(N87),.B(N1851));
AND2X1 AND2_354 (.Y(N2025),.A(N226),.B(N1852));
AND2X1 AND2_355 (.Y(N2026),.A(N97),.B(N1853));
AND2X1 AND2_356 (.Y(N2027),.A(N232),.B(N1854));
AND2X1 AND2_357 (.Y(N2028),.A(N107),.B(N1855));
AND2X1 AND2_358 (.Y(N2029),.A(N238),.B(N1856));
AND2X1 AND2_359 (.Y(N2030),.A(N116),.B(N1857));
AND2X1 AND2_360 (.Y(N2031),.A(N244),.B(N1858));
AND2X1 AND2_361 (.Y(N2032),.A(N283),.B(N1859));
AND2X1 AND2_362 (.Y(N2033),.A(N250),.B(N1860));
AND2X1 AND2_363 (.Y(N2034),.A(N294),.B(N1861));
AND2X1 AND2_364 (.Y(N2035),.A(N257),.B(N1862));
AND2X1 AND2_365 (.Y(N2036),.A(N303),.B(N1863));
AND2X1 AND2_366 (.Y(N2037),.A(N264),.B(N1864));
BUFX1 BUFF1_367 (.Y(N2038),.A(N1667));
INVX1 NOT1_368 (.Y(N2043),.A(N1667));
BUFX1 BUFF1_369 (.Y(N2052),.A(N1670));
INVX1 NOT1_370 (.Y(N2057),.A(N1670));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(N1197),.B(N1869));
AND2X1 AND_tmp61 (.Y(N2068),.A(N50),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(ttmp62),.A(N1197),.B(N1874));
AND2X1 AND_tmp63 (.Y(N2073),.A(N58),.B(ttmp62));
AND2X1 AND_tmp64 (.Y(ttmp64),.A(N1197),.B(N1879));
AND2X1 AND_tmp65 (.Y(N2078),.A(N68),.B(ttmp64));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(N1197),.B(N1884));
AND2X1 AND_tmp67 (.Y(N2083),.A(N77),.B(ttmp66));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(N1219),.B(N1889));
AND2X1 AND_tmp69 (.Y(N2088),.A(N87),.B(ttmp68));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(N1219),.B(N1894));
AND2X1 AND_tmp71 (.Y(N2093),.A(N97),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(ttmp72),.A(N1219),.B(N1899));
AND2X1 AND_tmp73 (.Y(N2098),.A(N107),.B(ttmp72));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(N1219),.B(N1904));
AND2X1 AND_tmp75 (.Y(N2103),.A(N116),.B(ttmp74));
INVX1 NOT1_379 (.Y(N2121),.A(N1562));
INVX1 NOT1_380 (.Y(N2122),.A(N1562));
INVX1 NOT1_381 (.Y(N2123),.A(N1562));
INVX1 NOT1_382 (.Y(N2124),.A(N1562));
INVX1 NOT1_383 (.Y(N2125),.A(N1562));
INVX1 NOT1_384 (.Y(N2126),.A(N1562));
INVX1 NOT1_385 (.Y(N2127),.A(N1562));
INVX1 NOT1_386 (.Y(N2128),.A(N1562));
NAND2X1 NAND2_387 (.Y(N2133),.A(N950),.B(N1939));
NAND2X1 NAND2_388 (.Y(N2134),.A(N1478),.B(N1941));
NAND2X1 NAND2_389 (.Y(N2135),.A(N1475),.B(N1942));
NAND2X1 NAND2_390 (.Y(N2136),.A(N1484),.B(N1943));
NAND2X1 NAND2_391 (.Y(N2137),.A(N1481),.B(N1944));
NAND2X1 NAND2_392 (.Y(N2138),.A(N1490),.B(N1945));
NAND2X1 NAND2_393 (.Y(N2139),.A(N1487),.B(N1946));
INVX1 NOT1_394 (.Y(N2141),.A(N1933));
INVX1 NOT1_395 (.Y(N2142),.A(N1936));
INVX1 NOT1_396 (.Y(N2143),.A(N1738));
AND2X1 AND2_397 (.Y(N2144),.A(N1738),.B(N1747));
INVX1 NOT1_398 (.Y(N2145),.A(N1747));
NAND2X1 NAND2_399 (.Y(N2146),.A(N1727),.B(N1960));
NAND2X1 NAND2_400 (.Y(N2147),.A(N1730),.B(N1961));
AND2X1 AND_tmp76 (.Y(ttmp76),.A(N665),.B(N58));
AND2X1 AND_tmp77 (.Y(ttmp77),.A(N1722),.B(ttmp76));
AND2X1 AND_tmp78 (.Y(N2148),.A(N1267),.B(ttmp77));
INVX1 NOT1_402 (.Y(N2149),.A(N1738));
AND2X1 AND2_403 (.Y(N2150),.A(N1738),.B(N1747));
INVX1 NOT1_404 (.Y(N2151),.A(N1747));
INVX1 NOT1_405 (.Y(N2152),.A(N1738));
INVX1 NOT1_406 (.Y(N2153),.A(N1747));
AND2X1 AND2_407 (.Y(N2154),.A(N1738),.B(N1747));
INVX1 NOT1_408 (.Y(N2155),.A(N1738));
INVX1 NOT1_409 (.Y(N2156),.A(N1747));
AND2X1 AND2_410 (.Y(N2157),.A(N1738),.B(N1747));
BUFX1 BUFF1_411 (.Y(N2158),.A(N1761));
BUFX1 BUFF1_412 (.Y(N2175),.A(N1761));
NAND2X1 NAND2_413 (.Y(N2178),.A(N1764),.B(N1981));
NAND2X1 NAND2_414 (.Y(N2179),.A(N1766),.B(N1982));
INVX1 NOT1_415 (.Y(N2180),.A(N1756));
AND2X1 AND2_416 (.Y(N2181),.A(N1756),.B(N1328));
INVX1 NOT1_417 (.Y(N2183),.A(N1756));
AND2X1 AND2_418 (.Y(N2184),.A(N1331),.B(N1756));
NAND2X1 NAND2_419 (.Y(N2185),.A(N1358),.B(N1812));
NAND2X1 NAND2_420 (.Y(N2188),.A(N1358),.B(N1809));
NAND2X1 NAND2_421 (.Y(N2191),.A(N1353),.B(N1812));
NAND2X1 NAND2_422 (.Y(N2194),.A(N1353),.B(N1809));
NAND2X1 NAND2_423 (.Y(N2197),.A(N1358),.B(N1806));
NAND2X1 NAND2_424 (.Y(N2200),.A(N1358),.B(N1803));
NAND2X1 NAND2_425 (.Y(N2203),.A(N1353),.B(N1806));
NAND2X1 NAND2_426 (.Y(N2206),.A(N1353),.B(N1803));
INVX1 NOT1_427 (.Y(N2209),.A(N1815));
INVX1 NOT1_428 (.Y(N2210),.A(N1818));
AND2X1 AND2_429 (.Y(N2211),.A(N1815),.B(N1818));
BUFX1 BUFF1_430 (.Y(N2212),.A(N1821));
BUFX1 BUFF1_431 (.Y(N2221),.A(N1821));
INVX1 NOT1_432 (.Y(N2230),.A(N1833));
INVX1 NOT1_433 (.Y(N2231),.A(N1833));
INVX1 NOT1_434 (.Y(N2232),.A(N1833));
INVX1 NOT1_435 (.Y(N2233),.A(N1833));
INVX1 NOT1_436 (.Y(N2234),.A(N1824));
INVX1 NOT1_437 (.Y(N2235),.A(N1824));
INVX1 NOT1_438 (.Y(N2236),.A(N1824));
INVX1 NOT1_439 (.Y(N2237),.A(N1824));
OR2X1 OR_tmp79 (.Y(ttmp79),.A(N1643),.B(N2023));
OR2X1 OR_tmp80 (.Y(N2238),.A(N2022),.B(ttmp79));
OR2X1 OR_tmp81 (.Y(ttmp81),.A(N1644),.B(N2025));
OR2X1 OR_tmp82 (.Y(N2239),.A(N2024),.B(ttmp81));
OR2X1 OR_tmp83 (.Y(ttmp83),.A(N1645),.B(N2027));
OR2X1 OR_tmp84 (.Y(N2240),.A(N2026),.B(ttmp83));
OR2X1 OR_tmp85 (.Y(ttmp85),.A(N1646),.B(N2029));
OR2X1 OR_tmp86 (.Y(N2241),.A(N2028),.B(ttmp85));
OR2X1 OR_tmp87 (.Y(ttmp87),.A(N1647),.B(N2031));
OR2X1 OR_tmp88 (.Y(N2242),.A(N2030),.B(ttmp87));
OR2X1 OR_tmp89 (.Y(ttmp89),.A(N1648),.B(N2033));
OR2X1 OR_tmp90 (.Y(N2243),.A(N2032),.B(ttmp89));
OR2X1 OR_tmp91 (.Y(ttmp91),.A(N1649),.B(N2035));
OR2X1 OR_tmp92 (.Y(N2244),.A(N2034),.B(ttmp91));
OR2X1 OR_tmp93 (.Y(ttmp93),.A(N1650),.B(N2037));
OR2X1 OR_tmp94 (.Y(N2245),.A(N2036),.B(ttmp93));
AND2X1 AND2_448 (.Y(N2270),.A(N1986),.B(N1673));
AND2X1 AND2_449 (.Y(N2277),.A(N1987),.B(N1675));
AND2X1 AND2_450 (.Y(N2282),.A(N1988),.B(N1676));
AND2X1 AND2_451 (.Y(N2287),.A(N1989),.B(N1677));
AND2X1 AND2_452 (.Y(N2294),.A(N1990),.B(N1679));
AND2X1 AND2_453 (.Y(N2299),.A(N1991),.B(N1680));
BUFX1 BUFF1_454 (.Y(N2304),.A(N1917));
AND2X1 AND2_455 (.Y(N2307),.A(N1930),.B(N350));
NAND2X1 NAND2_456 (.Y(N2310),.A(N1930),.B(N350));
BUFX1 BUFF1_457 (.Y(N2313),.A(N1715));
BUFX1 BUFF1_458 (.Y(N2316),.A(N1718));
BUFX1 BUFF1_459 (.Y(N2319),.A(N1715));
BUFX1 BUFF1_460 (.Y(N2322),.A(N1718));
NAND2X1 NAND2_461 (.Y(N2325),.A(N1940),.B(N2133));
NAND2X1 NAND2_462 (.Y(N2328),.A(N2134),.B(N2135));
NAND2X1 NAND2_463 (.Y(N2331),.A(N2136),.B(N2137));
NAND2X1 NAND2_464 (.Y(N2334),.A(N2138),.B(N2139));
NAND2X1 NAND2_465 (.Y(N2341),.A(N1936),.B(N2141));
NAND2X1 NAND2_466 (.Y(N2342),.A(N1933),.B(N2142));
AND2X1 AND2_467 (.Y(N2347),.A(N724),.B(N2144));
AND2X1 AND_tmp95 (.Y(ttmp95),.A(N699),.B(N1726));
AND2X1 AND_tmp96 (.Y(N2348),.A(N2146),.B(ttmp95));
AND2X1 AND2_469 (.Y(N2349),.A(N753),.B(N2147));
AND2X1 AND2_470 (.Y(N2350),.A(N2148),.B(N1273));
AND2X1 AND2_471 (.Y(N2351),.A(N736),.B(N2150));
AND2X1 AND2_472 (.Y(N2352),.A(N1735),.B(N2153));
AND2X1 AND2_473 (.Y(N2353),.A(N763),.B(N2154));
AND2X1 AND2_474 (.Y(N2354),.A(N1725),.B(N2156));
AND2X1 AND2_475 (.Y(N2355),.A(N749),.B(N2157));
INVX1 NOT1_476 (.Y(N2374),.A(N2178));
INVX1 NOT1_477 (.Y(N2375),.A(N2179));
AND2X1 AND2_478 (.Y(N2376),.A(N1520),.B(N2180));
AND2X1 AND2_479 (.Y(N2379),.A(N1721),.B(N2181));
AND2X1 AND2_480 (.Y(N2398),.A(N665),.B(N2211));
AND2X1 AND_tmp97 (.Y(ttmp97),.A(N226),.B(N1873));
AND2X1 AND_tmp98 (.Y(N2417),.A(N2057),.B(ttmp97));
AND2X1 AND_tmp99 (.Y(ttmp99),.A(N274),.B(N1306));
AND2X1 AND_tmp100 (.Y(N2418),.A(N2057),.B(ttmp99));
AND2X1 AND2_483 (.Y(N2419),.A(N2052),.B(N2238));
AND2X1 AND_tmp101 (.Y(ttmp101),.A(N232),.B(N1878));
AND2X1 AND_tmp102 (.Y(N2420),.A(N2057),.B(ttmp101));
AND2X1 AND_tmp103 (.Y(ttmp103),.A(N274),.B(N1306));
AND2X1 AND_tmp104 (.Y(N2421),.A(N2057),.B(ttmp103));
AND2X1 AND2_486 (.Y(N2422),.A(N2052),.B(N2239));
AND2X1 AND_tmp105 (.Y(ttmp105),.A(N238),.B(N1883));
AND2X1 AND_tmp106 (.Y(N2425),.A(N2057),.B(ttmp105));
AND2X1 AND_tmp107 (.Y(ttmp107),.A(N274),.B(N1306));
AND2X1 AND_tmp108 (.Y(N2426),.A(N2057),.B(ttmp107));
AND2X1 AND2_489 (.Y(N2427),.A(N2052),.B(N2240));
AND2X1 AND_tmp109 (.Y(ttmp109),.A(N244),.B(N1888));
AND2X1 AND_tmp110 (.Y(N2430),.A(N2057),.B(ttmp109));
AND2X1 AND_tmp111 (.Y(ttmp111),.A(N274),.B(N1306));
AND2X1 AND_tmp112 (.Y(N2431),.A(N2057),.B(ttmp111));
AND2X1 AND2_492 (.Y(N2432),.A(N2052),.B(N2241));
AND2X1 AND_tmp113 (.Y(ttmp113),.A(N250),.B(N1893));
AND2X1 AND_tmp114 (.Y(N2435),.A(N2043),.B(ttmp113));
AND2X1 AND_tmp115 (.Y(ttmp115),.A(N274),.B(N1322));
AND2X1 AND_tmp116 (.Y(N2436),.A(N2043),.B(ttmp115));
AND2X1 AND2_495 (.Y(N2437),.A(N2038),.B(N2242));
AND2X1 AND_tmp117 (.Y(ttmp117),.A(N257),.B(N1898));
AND2X1 AND_tmp118 (.Y(N2438),.A(N2043),.B(ttmp117));
AND2X1 AND_tmp119 (.Y(ttmp119),.A(N274),.B(N1315));
AND2X1 AND_tmp120 (.Y(N2439),.A(N2043),.B(ttmp119));
AND2X1 AND2_498 (.Y(N2440),.A(N2038),.B(N2243));
AND2X1 AND_tmp121 (.Y(ttmp121),.A(N264),.B(N1903));
AND2X1 AND_tmp122 (.Y(N2443),.A(N2043),.B(ttmp121));
AND2X1 AND_tmp123 (.Y(ttmp123),.A(N274),.B(N1315));
AND2X1 AND_tmp124 (.Y(N2444),.A(N2043),.B(ttmp123));
AND2X1 AND2_501 (.Y(N2445),.A(N2038),.B(N2244));
AND2X1 AND_tmp125 (.Y(ttmp125),.A(N270),.B(N1908));
AND2X1 AND_tmp126 (.Y(N2448),.A(N2043),.B(ttmp125));
AND2X1 AND_tmp127 (.Y(ttmp127),.A(N274),.B(N1315));
AND2X1 AND_tmp128 (.Y(N2449),.A(N2043),.B(ttmp127));
AND2X1 AND2_504 (.Y(N2450),.A(N2038),.B(N2245));
INVX1 NOT1_505 (.Y(N2467),.A(N2313));
INVX1 NOT1_506 (.Y(N2468),.A(N2316));
INVX1 NOT1_507 (.Y(N2469),.A(N2319));
INVX1 NOT1_508 (.Y(N2470),.A(N2322));
NAND2X1 NAND2_509 (.Y(N2471),.A(N2341),.B(N2342));
INVX1 NOT1_510 (.Y(N2474),.A(N2325));
INVX1 NOT1_511 (.Y(N2475),.A(N2328));
INVX1 NOT1_512 (.Y(N2476),.A(N2331));
INVX1 NOT1_513 (.Y(N2477),.A(N2334));
OR2X1 OR2_514 (.Y(N2478),.A(N2348),.B(N1729));
INVX1 NOT1_515 (.Y(N2481),.A(N2175));
AND2X1 AND2_516 (.Y(N2482),.A(N2175),.B(N1334));
AND2X1 AND2_517 (.Y(N2483),.A(N2349),.B(N2183));
AND2X1 AND2_518 (.Y(N2486),.A(N2374),.B(N1346));
AND2X1 AND2_519 (.Y(N2487),.A(N2375),.B(N1350));
BUFX1 BUFF1_520 (.Y(N2488),.A(N2185));
BUFX1 BUFF1_521 (.Y(N2497),.A(N2188));
BUFX1 BUFF1_522 (.Y(N2506),.A(N2191));
BUFX1 BUFF1_523 (.Y(N2515),.A(N2194));
BUFX1 BUFF1_524 (.Y(N2524),.A(N2197));
BUFX1 BUFF1_525 (.Y(N2533),.A(N2200));
BUFX1 BUFF1_526 (.Y(N2542),.A(N2203));
BUFX1 BUFF1_527 (.Y(N2551),.A(N2206));
BUFX1 BUFF1_528 (.Y(N2560),.A(N2185));
BUFX1 BUFF1_529 (.Y(N2569),.A(N2188));
BUFX1 BUFF1_530 (.Y(N2578),.A(N2191));
BUFX1 BUFF1_531 (.Y(N2587),.A(N2194));
BUFX1 BUFF1_532 (.Y(N2596),.A(N2197));
BUFX1 BUFF1_533 (.Y(N2605),.A(N2200));
BUFX1 BUFF1_534 (.Y(N2614),.A(N2203));
BUFX1 BUFF1_535 (.Y(N2623),.A(N2206));
INVX1 NOT1_536 (.Y(N2632),.A(N2212));
AND2X1 AND2_537 (.Y(N2633),.A(N2212),.B(N1833));
INVX1 NOT1_538 (.Y(N2634),.A(N2212));
AND2X1 AND2_539 (.Y(N2635),.A(N2212),.B(N1833));
INVX1 NOT1_540 (.Y(N2636),.A(N2212));
AND2X1 AND2_541 (.Y(N2637),.A(N2212),.B(N1833));
INVX1 NOT1_542 (.Y(N2638),.A(N2212));
AND2X1 AND2_543 (.Y(N2639),.A(N2212),.B(N1833));
INVX1 NOT1_544 (.Y(N2640),.A(N2221));
AND2X1 AND2_545 (.Y(N2641),.A(N2221),.B(N1824));
INVX1 NOT1_546 (.Y(N2642),.A(N2221));
AND2X1 AND2_547 (.Y(N2643),.A(N2221),.B(N1824));
INVX1 NOT1_548 (.Y(N2644),.A(N2221));
AND2X1 AND2_549 (.Y(N2645),.A(N2221),.B(N1824));
INVX1 NOT1_550 (.Y(N2646),.A(N2221));
AND2X1 AND2_551 (.Y(N2647),.A(N2221),.B(N1824));
OR2X1 OR_tmp129 (.Y(ttmp129),.A(N1870),.B(N2068));
OR2X1 OR_tmp130 (.Y(N2648),.A(N2270),.B(ttmp129));
OR2X1 OR_tmp131 (.Y(ttmp131),.A(N1870),.B(N2068));
NOR2X1 NOR_tmp132 (.Y(N2652),.A(N2270),.B(ttmp131));
OR2X1 OR_tmp133 (.Y(ttmp133),.A(N2418),.B(N2419));
OR2X1 OR_tmp134 (.Y(N2656),.A(N2417),.B(ttmp133));
OR2X1 OR_tmp135 (.Y(ttmp135),.A(N2421),.B(N2422));
OR2X1 OR_tmp136 (.Y(N2659),.A(N2420),.B(ttmp135));
OR2X1 OR_tmp137 (.Y(ttmp137),.A(N1880),.B(N2078));
OR2X1 OR_tmp138 (.Y(N2662),.A(N2277),.B(ttmp137));
OR2X1 OR_tmp139 (.Y(ttmp139),.A(N1880),.B(N2078));
NOR2X1 NOR_tmp140 (.Y(N2666),.A(N2277),.B(ttmp139));
OR2X1 OR_tmp141 (.Y(ttmp141),.A(N2426),.B(N2427));
OR2X1 OR_tmp142 (.Y(N2670),.A(N2425),.B(ttmp141));
OR2X1 OR_tmp143 (.Y(ttmp143),.A(N1885),.B(N2083));
OR2X1 OR_tmp144 (.Y(N2673),.A(N2282),.B(ttmp143));
OR2X1 OR_tmp145 (.Y(ttmp145),.A(N1885),.B(N2083));
NOR2X1 NOR_tmp146 (.Y(N2677),.A(N2282),.B(ttmp145));
OR2X1 OR_tmp147 (.Y(ttmp147),.A(N2431),.B(N2432));
OR2X1 OR_tmp148 (.Y(N2681),.A(N2430),.B(ttmp147));
OR2X1 OR_tmp149 (.Y(ttmp149),.A(N1890),.B(N2088));
OR2X1 OR_tmp150 (.Y(N2684),.A(N2287),.B(ttmp149));
OR2X1 OR_tmp151 (.Y(ttmp151),.A(N1890),.B(N2088));
NOR2X1 NOR_tmp152 (.Y(N2688),.A(N2287),.B(ttmp151));
OR2X1 OR_tmp153 (.Y(ttmp153),.A(N2436),.B(N2437));
OR2X1 OR_tmp154 (.Y(N2692),.A(N2435),.B(ttmp153));
OR2X1 OR_tmp155 (.Y(ttmp155),.A(N2439),.B(N2440));
OR2X1 OR_tmp156 (.Y(N2697),.A(N2438),.B(ttmp155));
OR2X1 OR_tmp157 (.Y(ttmp157),.A(N1900),.B(N2098));
OR2X1 OR_tmp158 (.Y(N2702),.A(N2294),.B(ttmp157));
OR2X1 OR_tmp159 (.Y(ttmp159),.A(N1900),.B(N2098));
NOR2X1 NOR_tmp160 (.Y(N2706),.A(N2294),.B(ttmp159));
OR2X1 OR_tmp161 (.Y(ttmp161),.A(N2444),.B(N2445));
OR2X1 OR_tmp162 (.Y(N2710),.A(N2443),.B(ttmp161));
OR2X1 OR_tmp163 (.Y(ttmp163),.A(N1905),.B(N2103));
OR2X1 OR_tmp164 (.Y(N2715),.A(N2299),.B(ttmp163));
OR2X1 OR_tmp165 (.Y(ttmp165),.A(N1905),.B(N2103));
NOR2X1 NOR_tmp166 (.Y(N2719),.A(N2299),.B(ttmp165));
OR2X1 OR_tmp167 (.Y(ttmp167),.A(N2449),.B(N2450));
OR2X1 OR_tmp168 (.Y(N2723),.A(N2448),.B(ttmp167));
INVX1 NOT1_572 (.Y(N2728),.A(N2304));
INVX1 NOT1_573 (.Y(N2729),.A(N2158));
AND2X1 AND2_574 (.Y(N2730),.A(N1562),.B(N2158));
INVX1 NOT1_575 (.Y(N2731),.A(N2158));
AND2X1 AND2_576 (.Y(N2732),.A(N1562),.B(N2158));
INVX1 NOT1_577 (.Y(N2733),.A(N2158));
AND2X1 AND2_578 (.Y(N2734),.A(N1562),.B(N2158));
INVX1 NOT1_579 (.Y(N2735),.A(N2158));
AND2X1 AND2_580 (.Y(N2736),.A(N1562),.B(N2158));
INVX1 NOT1_581 (.Y(N2737),.A(N2158));
AND2X1 AND2_582 (.Y(N2738),.A(N1562),.B(N2158));
INVX1 NOT1_583 (.Y(N2739),.A(N2158));
AND2X1 AND2_584 (.Y(N2740),.A(N1562),.B(N2158));
INVX1 NOT1_585 (.Y(N2741),.A(N2158));
AND2X1 AND2_586 (.Y(N2742),.A(N1562),.B(N2158));
INVX1 NOT1_587 (.Y(N2743),.A(N2158));
AND2X1 AND2_588 (.Y(N2744),.A(N1562),.B(N2158));
OR2X1 OR_tmp169 (.Y(ttmp169),.A(N1983),.B(N2379));
OR2X1 OR_tmp170 (.Y(N2745),.A(N2376),.B(ttmp169));
OR2X1 OR_tmp171 (.Y(ttmp171),.A(N1983),.B(N2379));
NOR2X1 NOR_tmp172 (.Y(N2746),.A(N2376),.B(ttmp171));
NAND2X1 NAND2_591 (.Y(N2748),.A(N2316),.B(N2467));
NAND2X1 NAND2_592 (.Y(N2749),.A(N2313),.B(N2468));
NAND2X1 NAND2_593 (.Y(N2750),.A(N2322),.B(N2469));
NAND2X1 NAND2_594 (.Y(N2751),.A(N2319),.B(N2470));
NAND2X1 NAND2_595 (.Y(N2754),.A(N2328),.B(N2474));
NAND2X1 NAND2_596 (.Y(N2755),.A(N2325),.B(N2475));
NAND2X1 NAND2_597 (.Y(N2756),.A(N2334),.B(N2476));
NAND2X1 NAND2_598 (.Y(N2757),.A(N2331),.B(N2477));
AND2X1 AND2_599 (.Y(N2758),.A(N1520),.B(N2481));
AND2X1 AND2_600 (.Y(N2761),.A(N1722),.B(N2482));
AND2X1 AND2_601 (.Y(N2764),.A(N2478),.B(N1770));
OR2X1 OR_tmp173 (.Y(ttmp173),.A(N1789),.B(N1790));
OR2X1 OR_tmp174 (.Y(N2768),.A(N2486),.B(ttmp173));
OR2X1 OR_tmp175 (.Y(ttmp175),.A(N1797),.B(N1798));
OR2X1 OR_tmp176 (.Y(N2769),.A(N2487),.B(ttmp175));
AND2X1 AND2_604 (.Y(N2898),.A(N665),.B(N2633));
AND2X1 AND2_605 (.Y(N2899),.A(N679),.B(N2635));
AND2X1 AND2_606 (.Y(N2900),.A(N686),.B(N2637));
AND2X1 AND2_607 (.Y(N2901),.A(N702),.B(N2639));
INVX1 NOT1_608 (.Y(N2962),.A(N2746));
NAND2X1 NAND2_609 (.Y(N2966),.A(N2748),.B(N2749));
NAND2X1 NAND2_610 (.Y(N2967),.A(N2750),.B(N2751));
BUFX1 BUFF1_611 (.Y(N2970),.A(N2471));
NAND2X1 NAND2_612 (.Y(N2973),.A(N2754),.B(N2755));
NAND2X1 NAND2_613 (.Y(N2977),.A(N2756),.B(N2757));
AND2X1 AND2_614 (.Y(N2980),.A(N2471),.B(N2143));
INVX1 NOT1_615 (.Y(N2984),.A(N2488));
INVX1 NOT1_616 (.Y(N2985),.A(N2497));
INVX1 NOT1_617 (.Y(N2986),.A(N2506));
INVX1 NOT1_618 (.Y(N2987),.A(N2515));
INVX1 NOT1_619 (.Y(N2988),.A(N2524));
INVX1 NOT1_620 (.Y(N2989),.A(N2533));
INVX1 NOT1_621 (.Y(N2990),.A(N2542));
INVX1 NOT1_622 (.Y(N2991),.A(N2551));
INVX1 NOT1_623 (.Y(N2992),.A(N2488));
INVX1 NOT1_624 (.Y(N2993),.A(N2497));
INVX1 NOT1_625 (.Y(N2994),.A(N2506));
INVX1 NOT1_626 (.Y(N2995),.A(N2515));
INVX1 NOT1_627 (.Y(N2996),.A(N2524));
INVX1 NOT1_628 (.Y(N2997),.A(N2533));
INVX1 NOT1_629 (.Y(N2998),.A(N2542));
INVX1 NOT1_630 (.Y(N2999),.A(N2551));
INVX1 NOT1_631 (.Y(N3000),.A(N2488));
INVX1 NOT1_632 (.Y(N3001),.A(N2497));
INVX1 NOT1_633 (.Y(N3002),.A(N2506));
INVX1 NOT1_634 (.Y(N3003),.A(N2515));
INVX1 NOT1_635 (.Y(N3004),.A(N2524));
INVX1 NOT1_636 (.Y(N3005),.A(N2533));
INVX1 NOT1_637 (.Y(N3006),.A(N2542));
INVX1 NOT1_638 (.Y(N3007),.A(N2551));
INVX1 NOT1_639 (.Y(N3008),.A(N2488));
INVX1 NOT1_640 (.Y(N3009),.A(N2497));
INVX1 NOT1_641 (.Y(N3010),.A(N2506));
INVX1 NOT1_642 (.Y(N3011),.A(N2515));
INVX1 NOT1_643 (.Y(N3012),.A(N2524));
INVX1 NOT1_644 (.Y(N3013),.A(N2533));
INVX1 NOT1_645 (.Y(N3014),.A(N2542));
INVX1 NOT1_646 (.Y(N3015),.A(N2551));
INVX1 NOT1_647 (.Y(N3016),.A(N2488));
INVX1 NOT1_648 (.Y(N3017),.A(N2497));
INVX1 NOT1_649 (.Y(N3018),.A(N2506));
INVX1 NOT1_650 (.Y(N3019),.A(N2515));
INVX1 NOT1_651 (.Y(N3020),.A(N2524));
INVX1 NOT1_652 (.Y(N3021),.A(N2533));
INVX1 NOT1_653 (.Y(N3022),.A(N2542));
INVX1 NOT1_654 (.Y(N3023),.A(N2551));
INVX1 NOT1_655 (.Y(N3024),.A(N2488));
INVX1 NOT1_656 (.Y(N3025),.A(N2497));
INVX1 NOT1_657 (.Y(N3026),.A(N2506));
INVX1 NOT1_658 (.Y(N3027),.A(N2515));
INVX1 NOT1_659 (.Y(N3028),.A(N2524));
INVX1 NOT1_660 (.Y(N3029),.A(N2533));
INVX1 NOT1_661 (.Y(N3030),.A(N2542));
INVX1 NOT1_662 (.Y(N3031),.A(N2551));
INVX1 NOT1_663 (.Y(N3032),.A(N2488));
INVX1 NOT1_664 (.Y(N3033),.A(N2497));
INVX1 NOT1_665 (.Y(N3034),.A(N2506));
INVX1 NOT1_666 (.Y(N3035),.A(N2515));
INVX1 NOT1_667 (.Y(N3036),.A(N2524));
INVX1 NOT1_668 (.Y(N3037),.A(N2533));
INVX1 NOT1_669 (.Y(N3038),.A(N2542));
INVX1 NOT1_670 (.Y(N3039),.A(N2551));
INVX1 NOT1_671 (.Y(N3040),.A(N2488));
INVX1 NOT1_672 (.Y(N3041),.A(N2497));
INVX1 NOT1_673 (.Y(N3042),.A(N2506));
INVX1 NOT1_674 (.Y(N3043),.A(N2515));
INVX1 NOT1_675 (.Y(N3044),.A(N2524));
INVX1 NOT1_676 (.Y(N3045),.A(N2533));
INVX1 NOT1_677 (.Y(N3046),.A(N2542));
INVX1 NOT1_678 (.Y(N3047),.A(N2551));
INVX1 NOT1_679 (.Y(N3048),.A(N2560));
INVX1 NOT1_680 (.Y(N3049),.A(N2569));
INVX1 NOT1_681 (.Y(N3050),.A(N2578));
INVX1 NOT1_682 (.Y(N3051),.A(N2587));
INVX1 NOT1_683 (.Y(N3052),.A(N2596));
INVX1 NOT1_684 (.Y(N3053),.A(N2605));
INVX1 NOT1_685 (.Y(N3054),.A(N2614));
INVX1 NOT1_686 (.Y(N3055),.A(N2623));
INVX1 NOT1_687 (.Y(N3056),.A(N2560));
INVX1 NOT1_688 (.Y(N3057),.A(N2569));
INVX1 NOT1_689 (.Y(N3058),.A(N2578));
INVX1 NOT1_690 (.Y(N3059),.A(N2587));
INVX1 NOT1_691 (.Y(N3060),.A(N2596));
INVX1 NOT1_692 (.Y(N3061),.A(N2605));
INVX1 NOT1_693 (.Y(N3062),.A(N2614));
INVX1 NOT1_694 (.Y(N3063),.A(N2623));
INVX1 NOT1_695 (.Y(N3064),.A(N2560));
INVX1 NOT1_696 (.Y(N3065),.A(N2569));
INVX1 NOT1_697 (.Y(N3066),.A(N2578));
INVX1 NOT1_698 (.Y(N3067),.A(N2587));
INVX1 NOT1_699 (.Y(N3068),.A(N2596));
INVX1 NOT1_700 (.Y(N3069),.A(N2605));
INVX1 NOT1_701 (.Y(N3070),.A(N2614));
INVX1 NOT1_702 (.Y(N3071),.A(N2623));
INVX1 NOT1_703 (.Y(N3072),.A(N2560));
INVX1 NOT1_704 (.Y(N3073),.A(N2569));
INVX1 NOT1_705 (.Y(N3074),.A(N2578));
INVX1 NOT1_706 (.Y(N3075),.A(N2587));
INVX1 NOT1_707 (.Y(N3076),.A(N2596));
INVX1 NOT1_708 (.Y(N3077),.A(N2605));
INVX1 NOT1_709 (.Y(N3078),.A(N2614));
INVX1 NOT1_710 (.Y(N3079),.A(N2623));
INVX1 NOT1_711 (.Y(N3080),.A(N2560));
INVX1 NOT1_712 (.Y(N3081),.A(N2569));
INVX1 NOT1_713 (.Y(N3082),.A(N2578));
INVX1 NOT1_714 (.Y(N3083),.A(N2587));
INVX1 NOT1_715 (.Y(N3084),.A(N2596));
INVX1 NOT1_716 (.Y(N3085),.A(N2605));
INVX1 NOT1_717 (.Y(N3086),.A(N2614));
INVX1 NOT1_718 (.Y(N3087),.A(N2623));
INVX1 NOT1_719 (.Y(N3088),.A(N2560));
INVX1 NOT1_720 (.Y(N3089),.A(N2569));
INVX1 NOT1_721 (.Y(N3090),.A(N2578));
INVX1 NOT1_722 (.Y(N3091),.A(N2587));
INVX1 NOT1_723 (.Y(N3092),.A(N2596));
INVX1 NOT1_724 (.Y(N3093),.A(N2605));
INVX1 NOT1_725 (.Y(N3094),.A(N2614));
INVX1 NOT1_726 (.Y(N3095),.A(N2623));
INVX1 NOT1_727 (.Y(N3096),.A(N2560));
INVX1 NOT1_728 (.Y(N3097),.A(N2569));
INVX1 NOT1_729 (.Y(N3098),.A(N2578));
INVX1 NOT1_730 (.Y(N3099),.A(N2587));
INVX1 NOT1_731 (.Y(N3100),.A(N2596));
INVX1 NOT1_732 (.Y(N3101),.A(N2605));
INVX1 NOT1_733 (.Y(N3102),.A(N2614));
INVX1 NOT1_734 (.Y(N3103),.A(N2623));
INVX1 NOT1_735 (.Y(N3104),.A(N2560));
INVX1 NOT1_736 (.Y(N3105),.A(N2569));
INVX1 NOT1_737 (.Y(N3106),.A(N2578));
INVX1 NOT1_738 (.Y(N3107),.A(N2587));
INVX1 NOT1_739 (.Y(N3108),.A(N2596));
INVX1 NOT1_740 (.Y(N3109),.A(N2605));
INVX1 NOT1_741 (.Y(N3110),.A(N2614));
INVX1 NOT1_742 (.Y(N3111),.A(N2623));
BUFX1 BUFF1_743 (.Y(N3112),.A(N2656));
INVX1 NOT1_744 (.Y(N3115),.A(N2656));
INVX1 NOT1_745 (.Y(N3118),.A(N2652));
AND2X1 AND2_746 (.Y(N3119),.A(N2768),.B(N1674));
BUFX1 BUFF1_747 (.Y(N3122),.A(N2659));
INVX1 NOT1_748 (.Y(N3125),.A(N2659));
BUFX1 BUFF1_749 (.Y(N3128),.A(N2670));
INVX1 NOT1_750 (.Y(N3131),.A(N2670));
INVX1 NOT1_751 (.Y(N3134),.A(N2666));
BUFX1 BUFF1_752 (.Y(N3135),.A(N2681));
INVX1 NOT1_753 (.Y(N3138),.A(N2681));
INVX1 NOT1_754 (.Y(N3141),.A(N2677));
BUFX1 BUFF1_755 (.Y(N3142),.A(N2692));
INVX1 NOT1_756 (.Y(N3145),.A(N2692));
INVX1 NOT1_757 (.Y(N3148),.A(N2688));
AND2X1 AND2_758 (.Y(N3149),.A(N2769),.B(N1678));
BUFX1 BUFF1_759 (.Y(N3152),.A(N2697));
INVX1 NOT1_760 (.Y(N3155),.A(N2697));
BUFX1 BUFF1_761 (.Y(N3158),.A(N2710));
INVX1 NOT1_762 (.Y(N3161),.A(N2710));
INVX1 NOT1_763 (.Y(N3164),.A(N2706));
BUFX1 BUFF1_764 (.Y(N3165),.A(N2723));
INVX1 NOT1_765 (.Y(N3168),.A(N2723));
INVX1 NOT1_766 (.Y(N3171),.A(N2719));
AND2X1 AND2_767 (.Y(N3172),.A(N1909),.B(N2648));
AND2X1 AND2_768 (.Y(N3175),.A(N1913),.B(N2662));
AND2X1 AND2_769 (.Y(N3178),.A(N1913),.B(N2673));
AND2X1 AND2_770 (.Y(N3181),.A(N1913),.B(N2684));
AND2X1 AND2_771 (.Y(N3184),.A(N1922),.B(N2702));
AND2X1 AND2_772 (.Y(N3187),.A(N1922),.B(N2715));
INVX1 NOT1_773 (.Y(N3190),.A(N2692));
INVX1 NOT1_774 (.Y(N3191),.A(N2697));
INVX1 NOT1_775 (.Y(N3192),.A(N2710));
INVX1 NOT1_776 (.Y(N3193),.A(N2723));
AND2X1 AND_tmp177 (.Y(ttmp177),.A(N2723),.B(N1459));
AND2X1 AND_tmp178 (.Y(ttmp178),.A(N2692),.B(ttmp177));
AND2X1 AND_tmp179 (.Y(ttmp179),.A(N2697),.B(ttmp178));
AND2X1 AND_tmp180 (.Y(N3194),.A(N2710),.B(ttmp179));
NAND2X1 NAND2_778 (.Y(N3195),.A(N2745),.B(N2962));
INVX1 NOT1_779 (.Y(N3196),.A(N2966));
OR2X1 OR_tmp181 (.Y(ttmp181),.A(N2145),.B(N2347));
OR2X1 OR_tmp182 (.Y(N3206),.A(N2980),.B(ttmp181));
AND2X1 AND2_781 (.Y(N3207),.A(N124),.B(N2984));
AND2X1 AND2_782 (.Y(N3208),.A(N159),.B(N2985));
AND2X1 AND2_783 (.Y(N3209),.A(N150),.B(N2986));
AND2X1 AND2_784 (.Y(N3210),.A(N143),.B(N2987));
AND2X1 AND2_785 (.Y(N3211),.A(N137),.B(N2988));
AND2X1 AND2_786 (.Y(N3212),.A(N132),.B(N2989));
AND2X1 AND2_787 (.Y(N3213),.A(N128),.B(N2990));
AND2X1 AND2_788 (.Y(N3214),.A(N125),.B(N2991));
AND2X1 AND2_789 (.Y(N3215),.A(N125),.B(N2992));
AND2X1 AND2_790 (.Y(N3216),.A(N655),.B(N2993));
AND2X1 AND2_791 (.Y(N3217),.A(N159),.B(N2994));
AND2X1 AND2_792 (.Y(N3218),.A(N150),.B(N2995));
AND2X1 AND2_793 (.Y(N3219),.A(N143),.B(N2996));
AND2X1 AND2_794 (.Y(N3220),.A(N137),.B(N2997));
AND2X1 AND2_795 (.Y(N3221),.A(N132),.B(N2998));
AND2X1 AND2_796 (.Y(N3222),.A(N128),.B(N2999));
AND2X1 AND2_797 (.Y(N3223),.A(N128),.B(N3000));
AND2X1 AND2_798 (.Y(N3224),.A(N670),.B(N3001));
AND2X1 AND2_799 (.Y(N3225),.A(N655),.B(N3002));
AND2X1 AND2_800 (.Y(N3226),.A(N159),.B(N3003));
AND2X1 AND2_801 (.Y(N3227),.A(N150),.B(N3004));
AND2X1 AND2_802 (.Y(N3228),.A(N143),.B(N3005));
AND2X1 AND2_803 (.Y(N3229),.A(N137),.B(N3006));
AND2X1 AND2_804 (.Y(N3230),.A(N132),.B(N3007));
AND2X1 AND2_805 (.Y(N3231),.A(N132),.B(N3008));
AND2X1 AND2_806 (.Y(N3232),.A(N690),.B(N3009));
AND2X1 AND2_807 (.Y(N3233),.A(N670),.B(N3010));
AND2X1 AND2_808 (.Y(N3234),.A(N655),.B(N3011));
AND2X1 AND2_809 (.Y(N3235),.A(N159),.B(N3012));
AND2X1 AND2_810 (.Y(N3236),.A(N150),.B(N3013));
AND2X1 AND2_811 (.Y(N3237),.A(N143),.B(N3014));
AND2X1 AND2_812 (.Y(N3238),.A(N137),.B(N3015));
AND2X1 AND2_813 (.Y(N3239),.A(N137),.B(N3016));
AND2X1 AND2_814 (.Y(N3240),.A(N706),.B(N3017));
AND2X1 AND2_815 (.Y(N3241),.A(N690),.B(N3018));
AND2X1 AND2_816 (.Y(N3242),.A(N670),.B(N3019));
AND2X1 AND2_817 (.Y(N3243),.A(N655),.B(N3020));
AND2X1 AND2_818 (.Y(N3244),.A(N159),.B(N3021));
AND2X1 AND2_819 (.Y(N3245),.A(N150),.B(N3022));
AND2X1 AND2_820 (.Y(N3246),.A(N143),.B(N3023));
AND2X1 AND2_821 (.Y(N3247),.A(N143),.B(N3024));
AND2X1 AND2_822 (.Y(N3248),.A(N715),.B(N3025));
AND2X1 AND2_823 (.Y(N3249),.A(N706),.B(N3026));
AND2X1 AND2_824 (.Y(N3250),.A(N690),.B(N3027));
AND2X1 AND2_825 (.Y(N3251),.A(N670),.B(N3028));
AND2X1 AND2_826 (.Y(N3252),.A(N655),.B(N3029));
AND2X1 AND2_827 (.Y(N3253),.A(N159),.B(N3030));
AND2X1 AND2_828 (.Y(N3254),.A(N150),.B(N3031));
AND2X1 AND2_829 (.Y(N3255),.A(N150),.B(N3032));
AND2X1 AND2_830 (.Y(N3256),.A(N727),.B(N3033));
AND2X1 AND2_831 (.Y(N3257),.A(N715),.B(N3034));
AND2X1 AND2_832 (.Y(N3258),.A(N706),.B(N3035));
AND2X1 AND2_833 (.Y(N3259),.A(N690),.B(N3036));
AND2X1 AND2_834 (.Y(N3260),.A(N670),.B(N3037));
AND2X1 AND2_835 (.Y(N3261),.A(N655),.B(N3038));
AND2X1 AND2_836 (.Y(N3262),.A(N159),.B(N3039));
AND2X1 AND2_837 (.Y(N3263),.A(N159),.B(N3040));
AND2X1 AND2_838 (.Y(N3264),.A(N740),.B(N3041));
AND2X1 AND2_839 (.Y(N3265),.A(N727),.B(N3042));
AND2X1 AND2_840 (.Y(N3266),.A(N715),.B(N3043));
AND2X1 AND2_841 (.Y(N3267),.A(N706),.B(N3044));
AND2X1 AND2_842 (.Y(N3268),.A(N690),.B(N3045));
AND2X1 AND2_843 (.Y(N3269),.A(N670),.B(N3046));
AND2X1 AND2_844 (.Y(N3270),.A(N655),.B(N3047));
AND2X1 AND2_845 (.Y(N3271),.A(N283),.B(N3048));
AND2X1 AND2_846 (.Y(N3272),.A(N670),.B(N3049));
AND2X1 AND2_847 (.Y(N3273),.A(N690),.B(N3050));
AND2X1 AND2_848 (.Y(N3274),.A(N706),.B(N3051));
AND2X1 AND2_849 (.Y(N3275),.A(N715),.B(N3052));
AND2X1 AND2_850 (.Y(N3276),.A(N727),.B(N3053));
AND2X1 AND2_851 (.Y(N3277),.A(N740),.B(N3054));
AND2X1 AND2_852 (.Y(N3278),.A(N753),.B(N3055));
AND2X1 AND2_853 (.Y(N3279),.A(N294),.B(N3056));
AND2X1 AND2_854 (.Y(N3280),.A(N690),.B(N3057));
AND2X1 AND2_855 (.Y(N3281),.A(N706),.B(N3058));
AND2X1 AND2_856 (.Y(N3282),.A(N715),.B(N3059));
AND2X1 AND2_857 (.Y(N3283),.A(N727),.B(N3060));
AND2X1 AND2_858 (.Y(N3284),.A(N740),.B(N3061));
AND2X1 AND2_859 (.Y(N3285),.A(N753),.B(N3062));
AND2X1 AND2_860 (.Y(N3286),.A(N283),.B(N3063));
AND2X1 AND2_861 (.Y(N3287),.A(N303),.B(N3064));
AND2X1 AND2_862 (.Y(N3288),.A(N706),.B(N3065));
AND2X1 AND2_863 (.Y(N3289),.A(N715),.B(N3066));
AND2X1 AND2_864 (.Y(N3290),.A(N727),.B(N3067));
AND2X1 AND2_865 (.Y(N3291),.A(N740),.B(N3068));
AND2X1 AND2_866 (.Y(N3292),.A(N753),.B(N3069));
AND2X1 AND2_867 (.Y(N3293),.A(N283),.B(N3070));
AND2X1 AND2_868 (.Y(N3294),.A(N294),.B(N3071));
AND2X1 AND2_869 (.Y(N3295),.A(N311),.B(N3072));
AND2X1 AND2_870 (.Y(N3296),.A(N715),.B(N3073));
AND2X1 AND2_871 (.Y(N3297),.A(N727),.B(N3074));
AND2X1 AND2_872 (.Y(N3298),.A(N740),.B(N3075));
AND2X1 AND2_873 (.Y(N3299),.A(N753),.B(N3076));
AND2X1 AND2_874 (.Y(N3300),.A(N283),.B(N3077));
AND2X1 AND2_875 (.Y(N3301),.A(N294),.B(N3078));
AND2X1 AND2_876 (.Y(N3302),.A(N303),.B(N3079));
AND2X1 AND2_877 (.Y(N3303),.A(N317),.B(N3080));
AND2X1 AND2_878 (.Y(N3304),.A(N727),.B(N3081));
AND2X1 AND2_879 (.Y(N3305),.A(N740),.B(N3082));
AND2X1 AND2_880 (.Y(N3306),.A(N753),.B(N3083));
AND2X1 AND2_881 (.Y(N3307),.A(N283),.B(N3084));
AND2X1 AND2_882 (.Y(N3308),.A(N294),.B(N3085));
AND2X1 AND2_883 (.Y(N3309),.A(N303),.B(N3086));
AND2X1 AND2_884 (.Y(N3310),.A(N311),.B(N3087));
AND2X1 AND2_885 (.Y(N3311),.A(N322),.B(N3088));
AND2X1 AND2_886 (.Y(N3312),.A(N740),.B(N3089));
AND2X1 AND2_887 (.Y(N3313),.A(N753),.B(N3090));
AND2X1 AND2_888 (.Y(N3314),.A(N283),.B(N3091));
AND2X1 AND2_889 (.Y(N3315),.A(N294),.B(N3092));
AND2X1 AND2_890 (.Y(N3316),.A(N303),.B(N3093));
AND2X1 AND2_891 (.Y(N3317),.A(N311),.B(N3094));
AND2X1 AND2_892 (.Y(N3318),.A(N317),.B(N3095));
AND2X1 AND2_893 (.Y(N3319),.A(N326),.B(N3096));
AND2X1 AND2_894 (.Y(N3320),.A(N753),.B(N3097));
AND2X1 AND2_895 (.Y(N3321),.A(N283),.B(N3098));
AND2X1 AND2_896 (.Y(N3322),.A(N294),.B(N3099));
AND2X1 AND2_897 (.Y(N3323),.A(N303),.B(N3100));
AND2X1 AND2_898 (.Y(N3324),.A(N311),.B(N3101));
AND2X1 AND2_899 (.Y(N3325),.A(N317),.B(N3102));
AND2X1 AND2_900 (.Y(N3326),.A(N322),.B(N3103));
AND2X1 AND2_901 (.Y(N3327),.A(N329),.B(N3104));
AND2X1 AND2_902 (.Y(N3328),.A(N283),.B(N3105));
AND2X1 AND2_903 (.Y(N3329),.A(N294),.B(N3106));
AND2X1 AND2_904 (.Y(N3330),.A(N303),.B(N3107));
AND2X1 AND2_905 (.Y(N3331),.A(N311),.B(N3108));
AND2X1 AND2_906 (.Y(N3332),.A(N317),.B(N3109));
AND2X1 AND2_907 (.Y(N3333),.A(N322),.B(N3110));
AND2X1 AND2_908 (.Y(N3334),.A(N326),.B(N3111));
AND2X1 AND_tmp183 (.Y(ttmp183),.A(N3193),.B(N917));
AND2X1 AND_tmp184 (.Y(ttmp184),.A(N3190),.B(ttmp183));
AND2X1 AND_tmp185 (.Y(ttmp185),.A(N3191),.B(ttmp184));
AND2X1 AND_tmp186 (.Y(N3383),.A(N3192),.B(ttmp185));
BUFX1 BUFF1_910 (.Y(N3384),.A(N2977));
AND2X1 AND2_911 (.Y(N3387),.A(N3196),.B(N1736));
AND2X1 AND2_912 (.Y(N3388),.A(N2977),.B(N2149));
AND2X1 AND2_913 (.Y(N3389),.A(N2973),.B(N1737));
OR2X1 OR_tmp187 (.Y(ttmp187),.A(N3213),.B(N3214));
OR2X1 OR_tmp188 (.Y(ttmp188),.A(N3207),.B(ttmp187));
OR2X1 OR_tmp189 (.Y(ttmp189),.A(N3208),.B(ttmp188));
OR2X1 OR_tmp190 (.Y(ttmp190),.A(N3209),.B(ttmp189));
OR2X1 OR_tmp191 (.Y(ttmp191),.A(N3210),.B(ttmp190));
OR2X1 OR_tmp192 (.Y(ttmp192),.A(N3211),.B(ttmp191));
NOR2X1 NOR_tmp193 (.Y(N3390),.A(N3212),.B(ttmp192));
OR2X1 OR_tmp194 (.Y(ttmp194),.A(N3221),.B(N3222));
OR2X1 OR_tmp195 (.Y(ttmp195),.A(N3215),.B(ttmp194));
OR2X1 OR_tmp196 (.Y(ttmp196),.A(N3216),.B(ttmp195));
OR2X1 OR_tmp197 (.Y(ttmp197),.A(N3217),.B(ttmp196));
OR2X1 OR_tmp198 (.Y(ttmp198),.A(N3218),.B(ttmp197));
OR2X1 OR_tmp199 (.Y(ttmp199),.A(N3219),.B(ttmp198));
NOR2X1 NOR_tmp200 (.Y(N3391),.A(N3220),.B(ttmp199));
OR2X1 OR_tmp201 (.Y(ttmp201),.A(N3229),.B(N3230));
OR2X1 OR_tmp202 (.Y(ttmp202),.A(N3223),.B(ttmp201));
OR2X1 OR_tmp203 (.Y(ttmp203),.A(N3224),.B(ttmp202));
OR2X1 OR_tmp204 (.Y(ttmp204),.A(N3225),.B(ttmp203));
OR2X1 OR_tmp205 (.Y(ttmp205),.A(N3226),.B(ttmp204));
OR2X1 OR_tmp206 (.Y(ttmp206),.A(N3227),.B(ttmp205));
NOR2X1 NOR_tmp207 (.Y(N3392),.A(N3228),.B(ttmp206));
OR2X1 OR_tmp208 (.Y(ttmp208),.A(N3237),.B(N3238));
OR2X1 OR_tmp209 (.Y(ttmp209),.A(N3231),.B(ttmp208));
OR2X1 OR_tmp210 (.Y(ttmp210),.A(N3232),.B(ttmp209));
OR2X1 OR_tmp211 (.Y(ttmp211),.A(N3233),.B(ttmp210));
OR2X1 OR_tmp212 (.Y(ttmp212),.A(N3234),.B(ttmp211));
OR2X1 OR_tmp213 (.Y(ttmp213),.A(N3235),.B(ttmp212));
NOR2X1 NOR_tmp214 (.Y(N3393),.A(N3236),.B(ttmp213));
OR2X1 OR_tmp215 (.Y(ttmp215),.A(N3245),.B(N3246));
OR2X1 OR_tmp216 (.Y(ttmp216),.A(N3239),.B(ttmp215));
OR2X1 OR_tmp217 (.Y(ttmp217),.A(N3240),.B(ttmp216));
OR2X1 OR_tmp218 (.Y(ttmp218),.A(N3241),.B(ttmp217));
OR2X1 OR_tmp219 (.Y(ttmp219),.A(N3242),.B(ttmp218));
OR2X1 OR_tmp220 (.Y(ttmp220),.A(N3243),.B(ttmp219));
NOR2X1 NOR_tmp221 (.Y(N3394),.A(N3244),.B(ttmp220));
OR2X1 OR_tmp222 (.Y(ttmp222),.A(N3253),.B(N3254));
OR2X1 OR_tmp223 (.Y(ttmp223),.A(N3247),.B(ttmp222));
OR2X1 OR_tmp224 (.Y(ttmp224),.A(N3248),.B(ttmp223));
OR2X1 OR_tmp225 (.Y(ttmp225),.A(N3249),.B(ttmp224));
OR2X1 OR_tmp226 (.Y(ttmp226),.A(N3250),.B(ttmp225));
OR2X1 OR_tmp227 (.Y(ttmp227),.A(N3251),.B(ttmp226));
NOR2X1 NOR_tmp228 (.Y(N3395),.A(N3252),.B(ttmp227));
OR2X1 OR_tmp229 (.Y(ttmp229),.A(N3261),.B(N3262));
OR2X1 OR_tmp230 (.Y(ttmp230),.A(N3255),.B(ttmp229));
OR2X1 OR_tmp231 (.Y(ttmp231),.A(N3256),.B(ttmp230));
OR2X1 OR_tmp232 (.Y(ttmp232),.A(N3257),.B(ttmp231));
OR2X1 OR_tmp233 (.Y(ttmp233),.A(N3258),.B(ttmp232));
OR2X1 OR_tmp234 (.Y(ttmp234),.A(N3259),.B(ttmp233));
NOR2X1 NOR_tmp235 (.Y(N3396),.A(N3260),.B(ttmp234));
OR2X1 OR_tmp236 (.Y(ttmp236),.A(N3269),.B(N3270));
OR2X1 OR_tmp237 (.Y(ttmp237),.A(N3263),.B(ttmp236));
OR2X1 OR_tmp238 (.Y(ttmp238),.A(N3264),.B(ttmp237));
OR2X1 OR_tmp239 (.Y(ttmp239),.A(N3265),.B(ttmp238));
OR2X1 OR_tmp240 (.Y(ttmp240),.A(N3266),.B(ttmp239));
OR2X1 OR_tmp241 (.Y(ttmp241),.A(N3267),.B(ttmp240));
NOR2X1 NOR_tmp242 (.Y(N3397),.A(N3268),.B(ttmp241));
OR2X1 OR_tmp243 (.Y(ttmp243),.A(N3277),.B(N3278));
OR2X1 OR_tmp244 (.Y(ttmp244),.A(N3271),.B(ttmp243));
OR2X1 OR_tmp245 (.Y(ttmp245),.A(N3272),.B(ttmp244));
OR2X1 OR_tmp246 (.Y(ttmp246),.A(N3273),.B(ttmp245));
OR2X1 OR_tmp247 (.Y(ttmp247),.A(N3274),.B(ttmp246));
OR2X1 OR_tmp248 (.Y(ttmp248),.A(N3275),.B(ttmp247));
NOR2X1 NOR_tmp249 (.Y(N3398),.A(N3276),.B(ttmp248));
OR2X1 OR_tmp250 (.Y(ttmp250),.A(N3285),.B(N3286));
OR2X1 OR_tmp251 (.Y(ttmp251),.A(N3279),.B(ttmp250));
OR2X1 OR_tmp252 (.Y(ttmp252),.A(N3280),.B(ttmp251));
OR2X1 OR_tmp253 (.Y(ttmp253),.A(N3281),.B(ttmp252));
OR2X1 OR_tmp254 (.Y(ttmp254),.A(N3282),.B(ttmp253));
OR2X1 OR_tmp255 (.Y(ttmp255),.A(N3283),.B(ttmp254));
NOR2X1 NOR_tmp256 (.Y(N3399),.A(N3284),.B(ttmp255));
OR2X1 OR_tmp257 (.Y(ttmp257),.A(N3293),.B(N3294));
OR2X1 OR_tmp258 (.Y(ttmp258),.A(N3287),.B(ttmp257));
OR2X1 OR_tmp259 (.Y(ttmp259),.A(N3288),.B(ttmp258));
OR2X1 OR_tmp260 (.Y(ttmp260),.A(N3289),.B(ttmp259));
OR2X1 OR_tmp261 (.Y(ttmp261),.A(N3290),.B(ttmp260));
OR2X1 OR_tmp262 (.Y(ttmp262),.A(N3291),.B(ttmp261));
NOR2X1 NOR_tmp263 (.Y(N3400),.A(N3292),.B(ttmp262));
OR2X1 OR_tmp264 (.Y(ttmp264),.A(N3301),.B(N3302));
OR2X1 OR_tmp265 (.Y(ttmp265),.A(N3295),.B(ttmp264));
OR2X1 OR_tmp266 (.Y(ttmp266),.A(N3296),.B(ttmp265));
OR2X1 OR_tmp267 (.Y(ttmp267),.A(N3297),.B(ttmp266));
OR2X1 OR_tmp268 (.Y(ttmp268),.A(N3298),.B(ttmp267));
OR2X1 OR_tmp269 (.Y(ttmp269),.A(N3299),.B(ttmp268));
NOR2X1 NOR_tmp270 (.Y(N3401),.A(N3300),.B(ttmp269));
OR2X1 OR_tmp271 (.Y(ttmp271),.A(N3309),.B(N3310));
OR2X1 OR_tmp272 (.Y(ttmp272),.A(N3303),.B(ttmp271));
OR2X1 OR_tmp273 (.Y(ttmp273),.A(N3304),.B(ttmp272));
OR2X1 OR_tmp274 (.Y(ttmp274),.A(N3305),.B(ttmp273));
OR2X1 OR_tmp275 (.Y(ttmp275),.A(N3306),.B(ttmp274));
OR2X1 OR_tmp276 (.Y(ttmp276),.A(N3307),.B(ttmp275));
NOR2X1 NOR_tmp277 (.Y(N3402),.A(N3308),.B(ttmp276));
OR2X1 OR_tmp278 (.Y(ttmp278),.A(N3317),.B(N3318));
OR2X1 OR_tmp279 (.Y(ttmp279),.A(N3311),.B(ttmp278));
OR2X1 OR_tmp280 (.Y(ttmp280),.A(N3312),.B(ttmp279));
OR2X1 OR_tmp281 (.Y(ttmp281),.A(N3313),.B(ttmp280));
OR2X1 OR_tmp282 (.Y(ttmp282),.A(N3314),.B(ttmp281));
OR2X1 OR_tmp283 (.Y(ttmp283),.A(N3315),.B(ttmp282));
NOR2X1 NOR_tmp284 (.Y(N3403),.A(N3316),.B(ttmp283));
OR2X1 OR_tmp285 (.Y(ttmp285),.A(N3325),.B(N3326));
OR2X1 OR_tmp286 (.Y(ttmp286),.A(N3319),.B(ttmp285));
OR2X1 OR_tmp287 (.Y(ttmp287),.A(N3320),.B(ttmp286));
OR2X1 OR_tmp288 (.Y(ttmp288),.A(N3321),.B(ttmp287));
OR2X1 OR_tmp289 (.Y(ttmp289),.A(N3322),.B(ttmp288));
OR2X1 OR_tmp290 (.Y(ttmp290),.A(N3323),.B(ttmp289));
NOR2X1 NOR_tmp291 (.Y(N3404),.A(N3324),.B(ttmp290));
OR2X1 OR_tmp292 (.Y(ttmp292),.A(N3333),.B(N3334));
OR2X1 OR_tmp293 (.Y(ttmp293),.A(N3327),.B(ttmp292));
OR2X1 OR_tmp294 (.Y(ttmp294),.A(N3328),.B(ttmp293));
OR2X1 OR_tmp295 (.Y(ttmp295),.A(N3329),.B(ttmp294));
OR2X1 OR_tmp296 (.Y(ttmp296),.A(N3330),.B(ttmp295));
OR2X1 OR_tmp297 (.Y(ttmp297),.A(N3331),.B(ttmp296));
NOR2X1 NOR_tmp298 (.Y(N3405),.A(N3332),.B(ttmp297));
AND2X1 AND2_930 (.Y(N3406),.A(N3206),.B(N2641));
AND2X1 AND_tmp299 (.Y(ttmp299),.A(N2648),.B(N3112));
AND2X1 AND_tmp300 (.Y(N3407),.A(N169),.B(ttmp299));
AND2X1 AND_tmp301 (.Y(ttmp301),.A(N2648),.B(N3115));
AND2X1 AND_tmp302 (.Y(N3410),.A(N179),.B(ttmp301));
AND2X1 AND_tmp303 (.Y(ttmp303),.A(N2652),.B(N3115));
AND2X1 AND_tmp304 (.Y(N3413),.A(N190),.B(ttmp303));
AND2X1 AND_tmp305 (.Y(ttmp305),.A(N2652),.B(N3112));
AND2X1 AND_tmp306 (.Y(N3414),.A(N200),.B(ttmp305));
OR2X1 OR_tmp307 (.Y(ttmp307),.A(N1875),.B(N2073));
OR2X1 OR_tmp308 (.Y(N3415),.A(N3119),.B(ttmp307));
OR2X1 OR_tmp309 (.Y(ttmp309),.A(N1875),.B(N2073));
NOR2X1 NOR_tmp310 (.Y(N3419),.A(N3119),.B(ttmp309));
AND2X1 AND_tmp311 (.Y(ttmp311),.A(N2662),.B(N3128));
AND2X1 AND_tmp312 (.Y(N3423),.A(N169),.B(ttmp311));
AND2X1 AND_tmp313 (.Y(ttmp313),.A(N2662),.B(N3131));
AND2X1 AND_tmp314 (.Y(N3426),.A(N179),.B(ttmp313));
AND2X1 AND_tmp315 (.Y(ttmp315),.A(N2666),.B(N3131));
AND2X1 AND_tmp316 (.Y(N3429),.A(N190),.B(ttmp315));
AND2X1 AND_tmp317 (.Y(ttmp317),.A(N2666),.B(N3128));
AND2X1 AND_tmp318 (.Y(N3430),.A(N200),.B(ttmp317));
AND2X1 AND_tmp319 (.Y(ttmp319),.A(N2673),.B(N3135));
AND2X1 AND_tmp320 (.Y(N3431),.A(N169),.B(ttmp319));
AND2X1 AND_tmp321 (.Y(ttmp321),.A(N2673),.B(N3138));
AND2X1 AND_tmp322 (.Y(N3434),.A(N179),.B(ttmp321));
AND2X1 AND_tmp323 (.Y(ttmp323),.A(N2677),.B(N3138));
AND2X1 AND_tmp324 (.Y(N3437),.A(N190),.B(ttmp323));
AND2X1 AND_tmp325 (.Y(ttmp325),.A(N2677),.B(N3135));
AND2X1 AND_tmp326 (.Y(N3438),.A(N200),.B(ttmp325));
AND2X1 AND_tmp327 (.Y(ttmp327),.A(N2684),.B(N3142));
AND2X1 AND_tmp328 (.Y(N3439),.A(N169),.B(ttmp327));
AND2X1 AND_tmp329 (.Y(ttmp329),.A(N2684),.B(N3145));
AND2X1 AND_tmp330 (.Y(N3442),.A(N179),.B(ttmp329));
AND2X1 AND_tmp331 (.Y(ttmp331),.A(N2688),.B(N3145));
AND2X1 AND_tmp332 (.Y(N3445),.A(N190),.B(ttmp331));
AND2X1 AND_tmp333 (.Y(ttmp333),.A(N2688),.B(N3142));
AND2X1 AND_tmp334 (.Y(N3446),.A(N200),.B(ttmp333));
OR2X1 OR_tmp335 (.Y(ttmp335),.A(N1895),.B(N2093));
OR2X1 OR_tmp336 (.Y(N3447),.A(N3149),.B(ttmp335));
OR2X1 OR_tmp337 (.Y(ttmp337),.A(N1895),.B(N2093));
NOR2X1 NOR_tmp338 (.Y(N3451),.A(N3149),.B(ttmp337));
AND2X1 AND_tmp339 (.Y(ttmp339),.A(N2702),.B(N3158));
AND2X1 AND_tmp340 (.Y(N3455),.A(N169),.B(ttmp339));
AND2X1 AND_tmp341 (.Y(ttmp341),.A(N2702),.B(N3161));
AND2X1 AND_tmp342 (.Y(N3458),.A(N179),.B(ttmp341));
AND2X1 AND_tmp343 (.Y(ttmp343),.A(N2706),.B(N3161));
AND2X1 AND_tmp344 (.Y(N3461),.A(N190),.B(ttmp343));
AND2X1 AND_tmp345 (.Y(ttmp345),.A(N2706),.B(N3158));
AND2X1 AND_tmp346 (.Y(N3462),.A(N200),.B(ttmp345));
AND2X1 AND_tmp347 (.Y(ttmp347),.A(N2715),.B(N3165));
AND2X1 AND_tmp348 (.Y(N3463),.A(N169),.B(ttmp347));
AND2X1 AND_tmp349 (.Y(ttmp349),.A(N2715),.B(N3168));
AND2X1 AND_tmp350 (.Y(N3466),.A(N179),.B(ttmp349));
AND2X1 AND_tmp351 (.Y(ttmp351),.A(N2719),.B(N3168));
AND2X1 AND_tmp352 (.Y(N3469),.A(N190),.B(ttmp351));
AND2X1 AND_tmp353 (.Y(ttmp353),.A(N2719),.B(N3165));
AND2X1 AND_tmp354 (.Y(N3470),.A(N200),.B(ttmp353));
OR2X1 OR2_959 (.Y(N3471),.A(N3194),.B(N3383));
BUFX1 BUFF1_960 (.Y(N3472),.A(N2967));
BUFX1 BUFF1_961 (.Y(N3475),.A(N2970));
BUFX1 BUFF1_962 (.Y(N3478),.A(N2967));
BUFX1 BUFF1_963 (.Y(N3481),.A(N2970));
BUFX1 BUFF1_964 (.Y(N3484),.A(N2973));
BUFX1 BUFF1_965 (.Y(N3487),.A(N2973));
BUFX1 BUFF1_966 (.Y(N3490),.A(N3172));
BUFX1 BUFF1_967 (.Y(N3493),.A(N3172));
BUFX1 BUFF1_968 (.Y(N3496),.A(N3175));
BUFX1 BUFF1_969 (.Y(N3499),.A(N3175));
BUFX1 BUFF1_970 (.Y(N3502),.A(N3178));
BUFX1 BUFF1_971 (.Y(N3505),.A(N3178));
BUFX1 BUFF1_972 (.Y(N3508),.A(N3181));
BUFX1 BUFF1_973 (.Y(N3511),.A(N3181));
BUFX1 BUFF1_974 (.Y(N3514),.A(N3184));
BUFX1 BUFF1_975 (.Y(N3517),.A(N3184));
BUFX1 BUFF1_976 (.Y(N3520),.A(N3187));
BUFX1 BUFF1_977 (.Y(N3523),.A(N3187));
NOR2X1 NOR2_978 (.Y(N3534),.A(N3387),.B(N2350));
OR2X1 OR_tmp355 (.Y(ttmp355),.A(N2151),.B(N2351));
OR2X1 OR_tmp356 (.Y(N3535),.A(N3388),.B(ttmp355));
NOR2X1 NOR2_980 (.Y(N3536),.A(N3389),.B(N1966));
AND2X1 AND2_981 (.Y(N3537),.A(N3390),.B(N2209));
AND2X1 AND2_982 (.Y(N3538),.A(N3398),.B(N2210));
AND2X1 AND2_983 (.Y(N3539),.A(N3391),.B(N1842));
AND2X1 AND2_984 (.Y(N3540),.A(N3399),.B(N1369));
AND2X1 AND2_985 (.Y(N3541),.A(N3392),.B(N1843));
AND2X1 AND2_986 (.Y(N3542),.A(N3400),.B(N1369));
AND2X1 AND2_987 (.Y(N3543),.A(N3393),.B(N1844));
AND2X1 AND2_988 (.Y(N3544),.A(N3401),.B(N1369));
AND2X1 AND2_989 (.Y(N3545),.A(N3394),.B(N1845));
AND2X1 AND2_990 (.Y(N3546),.A(N3402),.B(N1369));
AND2X1 AND2_991 (.Y(N3547),.A(N3395),.B(N1846));
AND2X1 AND2_992 (.Y(N3548),.A(N3403),.B(N1369));
AND2X1 AND2_993 (.Y(N3549),.A(N3396),.B(N1847));
AND2X1 AND2_994 (.Y(N3550),.A(N3404),.B(N1369));
AND2X1 AND2_995 (.Y(N3551),.A(N3397),.B(N1848));
AND2X1 AND2_996 (.Y(N3552),.A(N3405),.B(N1369));
OR2X1 OR_tmp357 (.Y(ttmp357),.A(N3414),.B(N3118));
OR2X1 OR_tmp358 (.Y(N3557),.A(N3413),.B(ttmp357));
OR2X1 OR_tmp359 (.Y(ttmp359),.A(N3430),.B(N3134));
OR2X1 OR_tmp360 (.Y(N3568),.A(N3429),.B(ttmp359));
OR2X1 OR_tmp361 (.Y(ttmp361),.A(N3438),.B(N3141));
OR2X1 OR_tmp362 (.Y(N3573),.A(N3437),.B(ttmp361));
OR2X1 OR_tmp363 (.Y(ttmp363),.A(N3446),.B(N3148));
OR2X1 OR_tmp364 (.Y(N3578),.A(N3445),.B(ttmp363));
OR2X1 OR_tmp365 (.Y(ttmp365),.A(N3462),.B(N3164));
OR2X1 OR_tmp366 (.Y(N3589),.A(N3461),.B(ttmp365));
OR2X1 OR_tmp367 (.Y(ttmp367),.A(N3470),.B(N3171));
OR2X1 OR_tmp368 (.Y(N3594),.A(N3469),.B(ttmp367));
AND2X1 AND2_1003 (.Y(N3605),.A(N3471),.B(N2728));
INVX1 NOT1_1004 (.Y(N3626),.A(N3478));
INVX1 NOT1_1005 (.Y(N3627),.A(N3481));
INVX1 NOT1_1006 (.Y(N3628),.A(N3487));
INVX1 NOT1_1007 (.Y(N3629),.A(N3484));
INVX1 NOT1_1008 (.Y(N3630),.A(N3472));
INVX1 NOT1_1009 (.Y(N3631),.A(N3475));
AND2X1 AND2_1010 (.Y(N3632),.A(N3536),.B(N2152));
AND2X1 AND2_1011 (.Y(N3633),.A(N3534),.B(N2155));
OR2X1 OR_tmp369 (.Y(ttmp369),.A(N3538),.B(N2398));
OR2X1 OR_tmp370 (.Y(N3634),.A(N3537),.B(ttmp369));
OR2X1 OR2_1013 (.Y(N3635),.A(N3539),.B(N3540));
OR2X1 OR2_1014 (.Y(N3636),.A(N3541),.B(N3542));
OR2X1 OR2_1015 (.Y(N3637),.A(N3543),.B(N3544));
OR2X1 OR2_1016 (.Y(N3638),.A(N3545),.B(N3546));
OR2X1 OR2_1017 (.Y(N3639),.A(N3547),.B(N3548));
OR2X1 OR2_1018 (.Y(N3640),.A(N3549),.B(N3550));
OR2X1 OR2_1019 (.Y(N3641),.A(N3551),.B(N3552));
AND2X1 AND2_1020 (.Y(N3642),.A(N3535),.B(N2643));
OR2X1 OR2_1021 (.Y(N3643),.A(N3407),.B(N3410));
NOR2X1 NOR2_1022 (.Y(N3644),.A(N3407),.B(N3410));
AND2X1 AND_tmp371 (.Y(ttmp371),.A(N3415),.B(N3122));
AND2X1 AND_tmp372 (.Y(N3645),.A(N169),.B(ttmp371));
AND2X1 AND_tmp373 (.Y(ttmp373),.A(N3415),.B(N3125));
AND2X1 AND_tmp374 (.Y(N3648),.A(N179),.B(ttmp373));
AND2X1 AND_tmp375 (.Y(ttmp375),.A(N3419),.B(N3125));
AND2X1 AND_tmp376 (.Y(N3651),.A(N190),.B(ttmp375));
AND2X1 AND_tmp377 (.Y(ttmp377),.A(N3419),.B(N3122));
AND2X1 AND_tmp378 (.Y(N3652),.A(N200),.B(ttmp377));
INVX1 NOT1_1027 (.Y(N3653),.A(N3419));
OR2X1 OR2_1028 (.Y(N3654),.A(N3423),.B(N3426));
NOR2X1 NOR2_1029 (.Y(N3657),.A(N3423),.B(N3426));
OR2X1 OR2_1030 (.Y(N3658),.A(N3431),.B(N3434));
NOR2X1 NOR2_1031 (.Y(N3661),.A(N3431),.B(N3434));
OR2X1 OR2_1032 (.Y(N3662),.A(N3439),.B(N3442));
NOR2X1 NOR2_1033 (.Y(N3663),.A(N3439),.B(N3442));
AND2X1 AND_tmp379 (.Y(ttmp379),.A(N3447),.B(N3152));
AND2X1 AND_tmp380 (.Y(N3664),.A(N169),.B(ttmp379));
AND2X1 AND_tmp381 (.Y(ttmp381),.A(N3447),.B(N3155));
AND2X1 AND_tmp382 (.Y(N3667),.A(N179),.B(ttmp381));
AND2X1 AND_tmp383 (.Y(ttmp383),.A(N3451),.B(N3155));
AND2X1 AND_tmp384 (.Y(N3670),.A(N190),.B(ttmp383));
AND2X1 AND_tmp385 (.Y(ttmp385),.A(N3451),.B(N3152));
AND2X1 AND_tmp386 (.Y(N3671),.A(N200),.B(ttmp385));
INVX1 NOT1_1038 (.Y(N3672),.A(N3451));
OR2X1 OR2_1039 (.Y(N3673),.A(N3455),.B(N3458));
NOR2X1 NOR2_1040 (.Y(N3676),.A(N3455),.B(N3458));
OR2X1 OR2_1041 (.Y(N3677),.A(N3463),.B(N3466));
NOR2X1 NOR2_1042 (.Y(N3680),.A(N3463),.B(N3466));
INVX1 NOT1_1043 (.Y(N3681),.A(N3493));
AND2X1 AND2_1044 (.Y(N3682),.A(N1909),.B(N3415));
INVX1 NOT1_1045 (.Y(N3685),.A(N3496));
INVX1 NOT1_1046 (.Y(N3686),.A(N3499));
INVX1 NOT1_1047 (.Y(N3687),.A(N3502));
INVX1 NOT1_1048 (.Y(N3688),.A(N3505));
INVX1 NOT1_1049 (.Y(N3689),.A(N3511));
AND2X1 AND2_1050 (.Y(N3690),.A(N1922),.B(N3447));
INVX1 NOT1_1051 (.Y(N3693),.A(N3517));
INVX1 NOT1_1052 (.Y(N3694),.A(N3520));
INVX1 NOT1_1053 (.Y(N3695),.A(N3523));
INVX1 NOT1_1054 (.Y(N3696),.A(N3514));
BUFX1 BUFF1_1055 (.Y(N3697),.A(N3384));
BUFX1 BUFF1_1056 (.Y(N3700),.A(N3384));
INVX1 NOT1_1057 (.Y(N3703),.A(N3490));
INVX1 NOT1_1058 (.Y(N3704),.A(N3508));
NAND2X1 NAND2_1059 (.Y(N3705),.A(N3475),.B(N3630));
NAND2X1 NAND2_1060 (.Y(N3706),.A(N3472),.B(N3631));
NAND2X1 NAND2_1061 (.Y(N3707),.A(N3481),.B(N3626));
NAND2X1 NAND2_1062 (.Y(N3708),.A(N3478),.B(N3627));
OR2X1 OR_tmp387 (.Y(ttmp387),.A(N2352),.B(N2353));
OR2X1 OR_tmp388 (.Y(N3711),.A(N3632),.B(ttmp387));
OR2X1 OR_tmp389 (.Y(ttmp389),.A(N2354),.B(N2355));
OR2X1 OR_tmp390 (.Y(N3712),.A(N3633),.B(ttmp389));
AND2X1 AND2_1065 (.Y(N3713),.A(N3634),.B(N2632));
AND2X1 AND2_1066 (.Y(N3714),.A(N3635),.B(N2634));
AND2X1 AND2_1067 (.Y(N3715),.A(N3636),.B(N2636));
AND2X1 AND2_1068 (.Y(N3716),.A(N3637),.B(N2638));
AND2X1 AND2_1069 (.Y(N3717),.A(N3638),.B(N2640));
AND2X1 AND2_1070 (.Y(N3718),.A(N3639),.B(N2642));
AND2X1 AND2_1071 (.Y(N3719),.A(N3640),.B(N2644));
AND2X1 AND2_1072 (.Y(N3720),.A(N3641),.B(N2646));
AND2X1 AND2_1073 (.Y(N3721),.A(N3644),.B(N3557));
OR2X1 OR_tmp391 (.Y(ttmp391),.A(N3652),.B(N3653));
OR2X1 OR_tmp392 (.Y(N3731),.A(N3651),.B(ttmp391));
AND2X1 AND2_1075 (.Y(N3734),.A(N3657),.B(N3568));
AND2X1 AND2_1076 (.Y(N3740),.A(N3661),.B(N3573));
AND2X1 AND2_1077 (.Y(N3743),.A(N3663),.B(N3578));
OR2X1 OR_tmp393 (.Y(ttmp393),.A(N3671),.B(N3672));
OR2X1 OR_tmp394 (.Y(N3753),.A(N3670),.B(ttmp393));
AND2X1 AND2_1079 (.Y(N3756),.A(N3676),.B(N3589));
AND2X1 AND2_1080 (.Y(N3762),.A(N3680),.B(N3594));
INVX1 NOT1_1081 (.Y(N3765),.A(N3643));
INVX1 NOT1_1082 (.Y(N3766),.A(N3662));
NAND2X1 NAND2_1083 (.Y(N3773),.A(N3705),.B(N3706));
NAND2X1 NAND2_1084 (.Y(N3774),.A(N3707),.B(N3708));
NAND2X1 NAND2_1085 (.Y(N3775),.A(N3700),.B(N3628));
INVX1 NOT1_1086 (.Y(N3776),.A(N3700));
NAND2X1 NAND2_1087 (.Y(N3777),.A(N3697),.B(N3629));
INVX1 NOT1_1088 (.Y(N3778),.A(N3697));
AND2X1 AND2_1089 (.Y(N3779),.A(N3712),.B(N2645));
AND2X1 AND2_1090 (.Y(N3780),.A(N3711),.B(N2647));
OR2X1 OR2_1091 (.Y(N3786),.A(N3645),.B(N3648));
NOR2X1 NOR2_1092 (.Y(N3789),.A(N3645),.B(N3648));
OR2X1 OR2_1093 (.Y(N3800),.A(N3664),.B(N3667));
NOR2X1 NOR2_1094 (.Y(N3803),.A(N3664),.B(N3667));
AND2X1 AND2_1095 (.Y(N3809),.A(N3654),.B(N1917));
AND2X1 AND2_1096 (.Y(N3812),.A(N3658),.B(N1917));
AND2X1 AND2_1097 (.Y(N3815),.A(N3673),.B(N1926));
AND2X1 AND2_1098 (.Y(N3818),.A(N3677),.B(N1926));
BUFX1 BUFF1_1099 (.Y(N3821),.A(N3682));
BUFX1 BUFF1_1100 (.Y(N3824),.A(N3682));
BUFX1 BUFF1_1101 (.Y(N3827),.A(N3690));
BUFX1 BUFF1_1102 (.Y(N3830),.A(N3690));
NAND2X1 NAND2_1103 (.Y(N3833),.A(N3773),.B(N3774));
NAND2X1 NAND2_1104 (.Y(N3834),.A(N3487),.B(N3776));
NAND2X1 NAND2_1105 (.Y(N3835),.A(N3484),.B(N3778));
AND2X1 AND2_1106 (.Y(N3838),.A(N3789),.B(N3731));
AND2X1 AND2_1107 (.Y(N3845),.A(N3803),.B(N3753));
BUFX1 BUFF1_1108 (.Y(N3850),.A(N3721));
BUFX1 BUFF1_1109 (.Y(N3855),.A(N3734));
BUFX1 BUFF1_1110 (.Y(N3858),.A(N3740));
BUFX1 BUFF1_1111 (.Y(N3861),.A(N3743));
BUFX1 BUFF1_1112 (.Y(N3865),.A(N3756));
BUFX1 BUFF1_1113 (.Y(N3868),.A(N3762));
NAND2X1 NAND2_1114 (.Y(N3884),.A(N3775),.B(N3834));
NAND2X1 NAND2_1115 (.Y(N3885),.A(N3777),.B(N3835));
NAND2X1 NAND2_1116 (.Y(N3894),.A(N3721),.B(N3786));
NAND2X1 NAND2_1117 (.Y(N3895),.A(N3743),.B(N3800));
INVX1 NOT1_1118 (.Y(N3898),.A(N3821));
INVX1 NOT1_1119 (.Y(N3899),.A(N3824));
INVX1 NOT1_1120 (.Y(N3906),.A(N3830));
INVX1 NOT1_1121 (.Y(N3911),.A(N3827));
AND2X1 AND2_1122 (.Y(N3912),.A(N3786),.B(N1912));
BUFX1 BUFF1_1123 (.Y(N3913),.A(N3812));
AND2X1 AND2_1124 (.Y(N3916),.A(N3800),.B(N1917));
BUFX1 BUFF1_1125 (.Y(N3917),.A(N3818));
INVX1 NOT1_1126 (.Y(N3920),.A(N3809));
BUFX1 BUFF1_1127 (.Y(N3921),.A(N3818));
INVX1 NOT1_1128 (.Y(N3924),.A(N3884));
INVX1 NOT1_1129 (.Y(N3925),.A(N3885));
AND2X1 AND_tmp395 (.Y(ttmp395),.A(N3734),.B(N3740));
AND2X1 AND_tmp396 (.Y(ttmp396),.A(N3721),.B(ttmp395));
AND2X1 AND_tmp397 (.Y(N3926),.A(N3838),.B(ttmp396));
AND2X1 AND_tmp398 (.Y(ttmp398),.A(N3838),.B(N3654));
NAND2X1 NAND_tmp399 (.Y(N3930),.A(N3721),.B(ttmp398));
AND2X1 AND_tmp400 (.Y(ttmp400),.A(N3734),.B(N3721));
AND2X1 AND_tmp401 (.Y(ttmp401),.A(N3658),.B(ttmp400));
NAND2X1 NAND_tmp402 (.Y(N3931),.A(N3838),.B(ttmp401));
AND2X1 AND_tmp403 (.Y(ttmp403),.A(N3756),.B(N3762));
AND2X1 AND_tmp404 (.Y(ttmp404),.A(N3743),.B(ttmp403));
AND2X1 AND_tmp405 (.Y(N3932),.A(N3845),.B(ttmp404));
AND2X1 AND_tmp406 (.Y(ttmp406),.A(N3845),.B(N3673));
NAND2X1 NAND_tmp407 (.Y(N3935),.A(N3743),.B(ttmp406));
AND2X1 AND_tmp408 (.Y(ttmp408),.A(N3756),.B(N3743));
AND2X1 AND_tmp409 (.Y(ttmp409),.A(N3677),.B(ttmp408));
NAND2X1 NAND_tmp410 (.Y(N3936),.A(N3845),.B(ttmp409));
BUFX1 BUFF1_1136 (.Y(N3937),.A(N3838));
BUFX1 BUFF1_1137 (.Y(N3940),.A(N3845));
INVX1 NOT1_1138 (.Y(N3947),.A(N3912));
INVX1 NOT1_1139 (.Y(N3948),.A(N3916));
BUFX1 BUFF1_1140 (.Y(N3950),.A(N3850));
BUFX1 BUFF1_1141 (.Y(N3953),.A(N3850));
BUFX1 BUFF1_1142 (.Y(N3956),.A(N3855));
BUFX1 BUFF1_1143 (.Y(N3959),.A(N3855));
BUFX1 BUFF1_1144 (.Y(N3962),.A(N3858));
BUFX1 BUFF1_1145 (.Y(N3965),.A(N3858));
BUFX1 BUFF1_1146 (.Y(N3968),.A(N3861));
BUFX1 BUFF1_1147 (.Y(N3971),.A(N3861));
BUFX1 BUFF1_1148 (.Y(N3974),.A(N3865));
BUFX1 BUFF1_1149 (.Y(N3977),.A(N3865));
BUFX1 BUFF1_1150 (.Y(N3980),.A(N3868));
BUFX1 BUFF1_1151 (.Y(N3983),.A(N3868));
NAND2X1 NAND2_1152 (.Y(N3987),.A(N3924),.B(N3925));
AND2X1 AND_tmp411 (.Y(ttmp411),.A(N3930),.B(N3931));
AND2X1 AND_tmp412 (.Y(ttmp412),.A(N3765),.B(ttmp411));
NAND2X1 NAND_tmp413 (.Y(N3992),.A(N3894),.B(ttmp412));
AND2X1 AND_tmp414 (.Y(ttmp414),.A(N3935),.B(N3936));
AND2X1 AND_tmp415 (.Y(ttmp415),.A(N3766),.B(ttmp414));
NAND2X1 NAND_tmp416 (.Y(N3996),.A(N3895),.B(ttmp415));
INVX1 NOT1_1155 (.Y(N4013),.A(N3921));
AND2X1 AND2_1156 (.Y(N4028),.A(N3932),.B(N3926));
NAND2X1 NAND2_1157 (.Y(N4029),.A(N3953),.B(N3681));
NAND2X1 NAND2_1158 (.Y(N4030),.A(N3959),.B(N3686));
NAND2X1 NAND2_1159 (.Y(N4031),.A(N3965),.B(N3688));
NAND2X1 NAND2_1160 (.Y(N4032),.A(N3971),.B(N3689));
NAND2X1 NAND2_1161 (.Y(N4033),.A(N3977),.B(N3693));
NAND2X1 NAND2_1162 (.Y(N4034),.A(N3983),.B(N3695));
BUFX1 BUFF1_1163 (.Y(N4035),.A(N3926));
INVX1 NOT1_1164 (.Y(N4042),.A(N3953));
INVX1 NOT1_1165 (.Y(N4043),.A(N3956));
NAND2X1 NAND2_1166 (.Y(N4044),.A(N3956),.B(N3685));
INVX1 NOT1_1167 (.Y(N4045),.A(N3959));
INVX1 NOT1_1168 (.Y(N4046),.A(N3962));
NAND2X1 NAND2_1169 (.Y(N4047),.A(N3962),.B(N3687));
INVX1 NOT1_1170 (.Y(N4048),.A(N3965));
INVX1 NOT1_1171 (.Y(N4049),.A(N3971));
INVX1 NOT1_1172 (.Y(N4050),.A(N3977));
INVX1 NOT1_1173 (.Y(N4051),.A(N3980));
NAND2X1 NAND2_1174 (.Y(N4052),.A(N3980),.B(N3694));
INVX1 NOT1_1175 (.Y(N4053),.A(N3983));
INVX1 NOT1_1176 (.Y(N4054),.A(N3974));
NAND2X1 NAND2_1177 (.Y(N4055),.A(N3974),.B(N3696));
AND2X1 AND2_1178 (.Y(N4056),.A(N3932),.B(N2304));
INVX1 NOT1_1179 (.Y(N4057),.A(N3950));
NAND2X1 NAND2_1180 (.Y(N4058),.A(N3950),.B(N3703));
BUFX1 BUFF1_1181 (.Y(N4059),.A(N3937));
BUFX1 BUFF1_1182 (.Y(N4062),.A(N3937));
INVX1 NOT1_1183 (.Y(N4065),.A(N3968));
NAND2X1 NAND2_1184 (.Y(N4066),.A(N3968),.B(N3704));
BUFX1 BUFF1_1185 (.Y(N4067),.A(N3940));
BUFX1 BUFF1_1186 (.Y(N4070),.A(N3940));
NAND2X1 NAND2_1187 (.Y(N4073),.A(N3926),.B(N3996));
INVX1 NOT1_1188 (.Y(N4074),.A(N3992));
NAND2X1 NAND2_1189 (.Y(N4075),.A(N3493),.B(N4042));
NAND2X1 NAND2_1190 (.Y(N4076),.A(N3499),.B(N4045));
NAND2X1 NAND2_1191 (.Y(N4077),.A(N3505),.B(N4048));
NAND2X1 NAND2_1192 (.Y(N4078),.A(N3511),.B(N4049));
NAND2X1 NAND2_1193 (.Y(N4079),.A(N3517),.B(N4050));
NAND2X1 NAND2_1194 (.Y(N4080),.A(N3523),.B(N4053));
NAND2X1 NAND2_1195 (.Y(N4085),.A(N3496),.B(N4043));
NAND2X1 NAND2_1196 (.Y(N4086),.A(N3502),.B(N4046));
NAND2X1 NAND2_1197 (.Y(N4088),.A(N3520),.B(N4051));
NAND2X1 NAND2_1198 (.Y(N4090),.A(N3514),.B(N4054));
AND2X1 AND2_1199 (.Y(N4091),.A(N3996),.B(N1926));
OR2X1 OR2_1200 (.Y(N4094),.A(N3605),.B(N4056));
NAND2X1 NAND2_1201 (.Y(N4098),.A(N3490),.B(N4057));
NAND2X1 NAND2_1202 (.Y(N4101),.A(N3508),.B(N4065));
AND2X1 AND2_1203 (.Y(N4104),.A(N4073),.B(N4074));
NAND2X1 NAND2_1204 (.Y(N4105),.A(N4075),.B(N4029));
NAND2X1 NAND2_1205 (.Y(N4106),.A(N4062),.B(N3899));
NAND2X1 NAND2_1206 (.Y(N4107),.A(N4076),.B(N4030));
NAND2X1 NAND2_1207 (.Y(N4108),.A(N4077),.B(N4031));
NAND2X1 NAND2_1208 (.Y(N4109),.A(N4078),.B(N4032));
NAND2X1 NAND2_1209 (.Y(N4110),.A(N4070),.B(N3906));
NAND2X1 NAND2_1210 (.Y(N4111),.A(N4079),.B(N4033));
NAND2X1 NAND2_1211 (.Y(N4112),.A(N4080),.B(N4034));
INVX1 NOT1_1212 (.Y(N4113),.A(N4059));
NAND2X1 NAND2_1213 (.Y(N4114),.A(N4059),.B(N3898));
INVX1 NOT1_1214 (.Y(N4115),.A(N4062));
NAND2X1 NAND2_1215 (.Y(N4116),.A(N4085),.B(N4044));
NAND2X1 NAND2_1216 (.Y(N4119),.A(N4086),.B(N4047));
INVX1 NOT1_1217 (.Y(N4122),.A(N4070));
NAND2X1 NAND2_1218 (.Y(N4123),.A(N4088),.B(N4052));
INVX1 NOT1_1219 (.Y(N4126),.A(N4067));
NAND2X1 NAND2_1220 (.Y(N4127),.A(N4067),.B(N3911));
NAND2X1 NAND2_1221 (.Y(N4128),.A(N4090),.B(N4055));
NAND2X1 NAND2_1222 (.Y(N4139),.A(N4098),.B(N4058));
NAND2X1 NAND2_1223 (.Y(N4142),.A(N4101),.B(N4066));
INVX1 NOT1_1224 (.Y(N4145),.A(N4104));
INVX1 NOT1_1225 (.Y(N4146),.A(N4105));
NAND2X1 NAND2_1226 (.Y(N4147),.A(N3824),.B(N4115));
INVX1 NOT1_1227 (.Y(N4148),.A(N4107));
INVX1 NOT1_1228 (.Y(N4149),.A(N4108));
INVX1 NOT1_1229 (.Y(N4150),.A(N4109));
NAND2X1 NAND2_1230 (.Y(N4151),.A(N3830),.B(N4122));
INVX1 NOT1_1231 (.Y(N4152),.A(N4111));
INVX1 NOT1_1232 (.Y(N4153),.A(N4112));
NAND2X1 NAND2_1233 (.Y(N4154),.A(N3821),.B(N4113));
NAND2X1 NAND2_1234 (.Y(N4161),.A(N3827),.B(N4126));
BUFX1 BUFF1_1235 (.Y(N4167),.A(N4091));
BUFX1 BUFF1_1236 (.Y(N4174),.A(N4094));
BUFX1 BUFF1_1237 (.Y(N4182),.A(N4091));
AND2X1 AND2_1238 (.Y(N4186),.A(N330),.B(N4094));
AND2X1 AND2_1239 (.Y(N4189),.A(N4146),.B(N2230));
NAND2X1 NAND2_1240 (.Y(N4190),.A(N4147),.B(N4106));
AND2X1 AND2_1241 (.Y(N4191),.A(N4148),.B(N2232));
AND2X1 AND2_1242 (.Y(N4192),.A(N4149),.B(N2233));
AND2X1 AND2_1243 (.Y(N4193),.A(N4150),.B(N2234));
NAND2X1 NAND2_1244 (.Y(N4194),.A(N4151),.B(N4110));
AND2X1 AND2_1245 (.Y(N4195),.A(N4152),.B(N2236));
AND2X1 AND2_1246 (.Y(N4196),.A(N4153),.B(N2237));
NAND2X1 NAND2_1247 (.Y(N4197),.A(N4154),.B(N4114));
BUFX1 BUFF1_1248 (.Y(N4200),.A(N4116));
BUFX1 BUFF1_1249 (.Y(N4203),.A(N4116));
BUFX1 BUFF1_1250 (.Y(N4209),.A(N4119));
BUFX1 BUFF1_1251 (.Y(N4213),.A(N4119));
NAND2X1 NAND2_1252 (.Y(N4218),.A(N4161),.B(N4127));
BUFX1 BUFF1_1253 (.Y(N4223),.A(N4123));
AND2X1 AND2_1254 (.Y(N4238),.A(N4128),.B(N3917));
INVX1 NOT1_1255 (.Y(N4239),.A(N4139));
INVX1 NOT1_1256 (.Y(N4241),.A(N4142));
AND2X1 AND2_1257 (.Y(N4242),.A(N330),.B(N4123));
BUFX1 BUFF1_1258 (.Y(N4247),.A(N4128));
OR2X1 OR_tmp417 (.Y(ttmp417),.A(N4189),.B(N2898));
NOR2X1 NOR_tmp418 (.Y(N4251),.A(N3713),.B(ttmp417));
INVX1 NOT1_1260 (.Y(N4252),.A(N4190));
OR2X1 OR_tmp419 (.Y(ttmp419),.A(N4191),.B(N2900));
NOR2X1 NOR_tmp420 (.Y(N4253),.A(N3715),.B(ttmp419));
OR2X1 OR_tmp421 (.Y(ttmp421),.A(N4192),.B(N2901));
NOR2X1 NOR_tmp422 (.Y(N4254),.A(N3716),.B(ttmp421));
OR2X1 OR_tmp423 (.Y(ttmp423),.A(N4193),.B(N3406));
NOR2X1 NOR_tmp424 (.Y(N4255),.A(N3717),.B(ttmp423));
INVX1 NOT1_1264 (.Y(N4256),.A(N4194));
OR2X1 OR_tmp425 (.Y(ttmp425),.A(N4195),.B(N3779));
NOR2X1 NOR_tmp426 (.Y(N4257),.A(N3719),.B(ttmp425));
OR2X1 OR_tmp427 (.Y(ttmp427),.A(N4196),.B(N3780));
NOR2X1 NOR_tmp428 (.Y(N4258),.A(N3720),.B(ttmp427));
AND2X1 AND2_1267 (.Y(N4283),.A(N4167),.B(N4035));
AND2X1 AND2_1268 (.Y(N4284),.A(N4174),.B(N4035));
OR2X1 OR2_1269 (.Y(N4287),.A(N3815),.B(N4238));
INVX1 NOT1_1270 (.Y(N4291),.A(N4186));
INVX1 NOT1_1271 (.Y(N4295),.A(N4167));
BUFX1 BUFF1_1272 (.Y(N4296),.A(N4167));
INVX1 NOT1_1273 (.Y(N4299),.A(N4182));
AND2X1 AND2_1274 (.Y(N4303),.A(N4252),.B(N2231));
AND2X1 AND2_1275 (.Y(N4304),.A(N4256),.B(N2235));
BUFX1 BUFF1_1276 (.Y(N4305),.A(N4197));
OR2X1 OR2_1277 (.Y(N4310),.A(N3992),.B(N4283));
AND2X1 AND_tmp429 (.Y(ttmp429),.A(N4213),.B(N4203));
AND2X1 AND_tmp430 (.Y(N4316),.A(N4174),.B(ttmp429));
AND2X1 AND2_1279 (.Y(N4317),.A(N4174),.B(N4209));
AND2X1 AND_tmp431 (.Y(ttmp431),.A(N4128),.B(N4218));
AND2X1 AND_tmp432 (.Y(N4318),.A(N4223),.B(ttmp431));
AND2X1 AND2_1281 (.Y(N4319),.A(N4223),.B(N4128));
AND2X1 AND2_1282 (.Y(N4322),.A(N4167),.B(N4209));
NAND2X1 NAND2_1283 (.Y(N4325),.A(N4203),.B(N3913));
AND2X1 AND_tmp433 (.Y(ttmp433),.A(N4213),.B(N4167));
NAND2X1 NAND_tmp434 (.Y(N4326),.A(N4203),.B(ttmp433));
NAND2X1 NAND2_1285 (.Y(N4327),.A(N4218),.B(N3815));
AND2X1 AND_tmp435 (.Y(ttmp435),.A(N4128),.B(N3917));
NAND2X1 NAND_tmp436 (.Y(N4328),.A(N4218),.B(ttmp435));
NAND2X1 NAND2_1287 (.Y(N4329),.A(N4247),.B(N4013));
INVX1 NOT1_1288 (.Y(N4330),.A(N4247));
AND2X1 AND_tmp437 (.Y(ttmp437),.A(N4094),.B(N4295));
AND2X1 AND_tmp438 (.Y(N4331),.A(N330),.B(ttmp437));
AND2X1 AND2_1290 (.Y(N4335),.A(N4251),.B(N2730));
AND2X1 AND2_1291 (.Y(N4338),.A(N4253),.B(N2734));
AND2X1 AND2_1292 (.Y(N4341),.A(N4254),.B(N2736));
AND2X1 AND2_1293 (.Y(N4344),.A(N4255),.B(N2738));
AND2X1 AND2_1294 (.Y(N4347),.A(N4257),.B(N2742));
AND2X1 AND2_1295 (.Y(N4350),.A(N4258),.B(N2744));
BUFX1 BUFF1_1296 (.Y(N4353),.A(N4197));
BUFX1 BUFF1_1297 (.Y(N4356),.A(N4203));
BUFX1 BUFF1_1298 (.Y(N4359),.A(N4209));
BUFX1 BUFF1_1299 (.Y(N4362),.A(N4218));
BUFX1 BUFF1_1300 (.Y(N4365),.A(N4242));
BUFX1 BUFF1_1301 (.Y(N4368),.A(N4242));
AND2X1 AND2_1302 (.Y(N4371),.A(N4223),.B(N4223));
OR2X1 OR_tmp439 (.Y(ttmp439),.A(N4303),.B(N2899));
NOR2X1 NOR_tmp440 (.Y(N4376),.A(N3714),.B(ttmp439));
OR2X1 OR_tmp441 (.Y(ttmp441),.A(N4304),.B(N3642));
NOR2X1 NOR_tmp442 (.Y(N4377),.A(N3718),.B(ttmp441));
AND2X1 AND2_1305 (.Y(N4387),.A(N330),.B(N4317));
AND2X1 AND2_1306 (.Y(N4390),.A(N330),.B(N4318));
NAND2X1 NAND2_1307 (.Y(N4393),.A(N3921),.B(N4330));
BUFX1 BUFF1_1308 (.Y(N4398),.A(N4287));
BUFX1 BUFF1_1309 (.Y(N4413),.A(N4284));
AND2X1 AND_tmp443 (.Y(ttmp443),.A(N4325),.B(N4326));
NAND2X1 NAND_tmp444 (.Y(N4416),.A(N3920),.B(ttmp443));
OR2X1 OR2_1311 (.Y(N4421),.A(N3812),.B(N4322));
AND2X1 AND_tmp445 (.Y(ttmp445),.A(N4327),.B(N4328));
NAND2X1 NAND_tmp446 (.Y(N4427),.A(N3948),.B(ttmp445));
BUFX1 BUFF1_1313 (.Y(N4430),.A(N4287));
AND2X1 AND2_1314 (.Y(N4435),.A(N330),.B(N4316));
OR2X1 OR2_1315 (.Y(N4442),.A(N4331),.B(N4296));
AND2X1 AND_tmp447 (.Y(ttmp447),.A(N4203),.B(N4213));
AND2X1 AND_tmp448 (.Y(ttmp448),.A(N4174),.B(ttmp447));
AND2X1 AND_tmp449 (.Y(N4443),.A(N4305),.B(ttmp448));
NAND2X1 NAND2_1317 (.Y(N4446),.A(N4305),.B(N3809));
AND2X1 AND_tmp450 (.Y(ttmp450),.A(N4200),.B(N3913));
NAND2X1 NAND_tmp451 (.Y(N4447),.A(N4305),.B(ttmp450));
AND2X1 AND_tmp452 (.Y(ttmp452),.A(N4213),.B(N4167));
AND2X1 AND_tmp453 (.Y(ttmp453),.A(N4305),.B(ttmp452));
NAND2X1 NAND_tmp454 (.Y(N4448),.A(N4200),.B(ttmp453));
INVX1 NOT1_1320 (.Y(N4452),.A(N4356));
NAND2X1 NAND2_1321 (.Y(N4458),.A(N4329),.B(N4393));
INVX1 NOT1_1322 (.Y(N4461),.A(N4365));
INVX1 NOT1_1323 (.Y(N4462),.A(N4368));
NAND2X1 NAND2_1324 (.Y(N4463),.A(N4371),.B(N1460));
INVX1 NOT1_1325 (.Y(N4464),.A(N4371));
BUFX1 BUFF1_1326 (.Y(N4465),.A(N4310));
NOR2X1 NOR2_1327 (.Y(N4468),.A(N4331),.B(N4296));
AND2X1 AND2_1328 (.Y(N4472),.A(N4376),.B(N2732));
AND2X1 AND2_1329 (.Y(N4475),.A(N4377),.B(N2740));
BUFX1 BUFF1_1330 (.Y(N4479),.A(N4310));
INVX1 NOT1_1331 (.Y(N4484),.A(N4353));
INVX1 NOT1_1332 (.Y(N4486),.A(N4359));
NAND2X1 NAND2_1333 (.Y(N4487),.A(N4359),.B(N4299));
INVX1 NOT1_1334 (.Y(N4491),.A(N4362));
AND2X1 AND2_1335 (.Y(N4493),.A(N330),.B(N4319));
INVX1 NOT1_1336 (.Y(N4496),.A(N4398));
AND2X1 AND2_1337 (.Y(N4497),.A(N4287),.B(N4398));
AND2X1 AND2_1338 (.Y(N4498),.A(N4442),.B(N1769));
AND2X1 AND_tmp455 (.Y(ttmp455),.A(N4447),.B(N4448));
AND2X1 AND_tmp456 (.Y(ttmp456),.A(N3947),.B(ttmp455));
NAND2X1 NAND_tmp457 (.Y(N4503),.A(N4446),.B(ttmp456));
INVX1 NOT1_1340 (.Y(N4506),.A(N4413));
INVX1 NOT1_1341 (.Y(N4507),.A(N4435));
INVX1 NOT1_1342 (.Y(N4508),.A(N4421));
NAND2X1 NAND2_1343 (.Y(N4509),.A(N4421),.B(N4452));
INVX1 NOT1_1344 (.Y(N4510),.A(N4427));
NAND2X1 NAND2_1345 (.Y(N4511),.A(N4427),.B(N4241));
NAND2X1 NAND2_1346 (.Y(N4515),.A(N965),.B(N4464));
INVX1 NOT1_1347 (.Y(N4526),.A(N4416));
NAND2X1 NAND2_1348 (.Y(N4527),.A(N4416),.B(N4484));
NAND2X1 NAND2_1349 (.Y(N4528),.A(N4182),.B(N4486));
INVX1 NOT1_1350 (.Y(N4529),.A(N4430));
NAND2X1 NAND2_1351 (.Y(N4530),.A(N4430),.B(N4491));
BUFX1 BUFF1_1352 (.Y(N4531),.A(N4387));
BUFX1 BUFF1_1353 (.Y(N4534),.A(N4387));
BUFX1 BUFF1_1354 (.Y(N4537),.A(N4390));
BUFX1 BUFF1_1355 (.Y(N4540),.A(N4390));
AND2X1 AND_tmp458 (.Y(ttmp458),.A(N4319),.B(N4496));
AND2X1 AND_tmp459 (.Y(N4545),.A(N330),.B(ttmp458));
AND2X1 AND2_1357 (.Y(N4549),.A(N330),.B(N4443));
NAND2X1 NAND2_1358 (.Y(N4552),.A(N4356),.B(N4508));
NAND2X1 NAND2_1359 (.Y(N4555),.A(N4142),.B(N4510));
INVX1 NOT1_1360 (.Y(N4558),.A(N4493));
NAND2X1 NAND2_1361 (.Y(N4559),.A(N4463),.B(N4515));
INVX1 NOT1_1362 (.Y(N4562),.A(N4465));
AND2X1 AND2_1363 (.Y(N4563),.A(N4310),.B(N4465));
BUFX1 BUFF1_1364 (.Y(N4564),.A(N4468));
INVX1 NOT1_1365 (.Y(N4568),.A(N4479));
BUFX1 BUFF1_1366 (.Y(N4569),.A(N4443));
NAND2X1 NAND2_1367 (.Y(N4572),.A(N4353),.B(N4526));
NAND2X1 NAND2_1368 (.Y(N4573),.A(N4362),.B(N4529));
NAND2X1 NAND2_1369 (.Y(N4576),.A(N4487),.B(N4528));
BUFX1 BUFF1_1370 (.Y(N4581),.A(N4458));
BUFX1 BUFF1_1371 (.Y(N4584),.A(N4458));
OR2X1 OR_tmp460 (.Y(ttmp460),.A(N4498),.B(N2761));
OR2X1 OR_tmp461 (.Y(N4587),.A(N2758),.B(ttmp460));
OR2X1 OR_tmp462 (.Y(ttmp462),.A(N4498),.B(N2761));
NOR2X1 NOR_tmp463 (.Y(N4588),.A(N2758),.B(ttmp462));
OR2X1 OR2_1374 (.Y(N4589),.A(N4545),.B(N4497));
NAND2X1 NAND2_1375 (.Y(N4593),.A(N4552),.B(N4509));
INVX1 NOT1_1376 (.Y(N4596),.A(N4531));
INVX1 NOT1_1377 (.Y(N4597),.A(N4534));
NAND2X1 NAND2_1378 (.Y(N4599),.A(N4555),.B(N4511));
INVX1 NOT1_1379 (.Y(N4602),.A(N4537));
INVX1 NOT1_1380 (.Y(N4603),.A(N4540));
AND2X1 AND_tmp464 (.Y(ttmp464),.A(N4284),.B(N4562));
AND2X1 AND_tmp465 (.Y(N4608),.A(N330),.B(ttmp464));
BUFX1 BUFF1_1382 (.Y(N4613),.A(N4503));
BUFX1 BUFF1_1383 (.Y(N4616),.A(N4503));
NAND2X1 NAND2_1384 (.Y(N4619),.A(N4572),.B(N4527));
NAND2X1 NAND2_1385 (.Y(N4623),.A(N4573),.B(N4530));
INVX1 NOT1_1386 (.Y(N4628),.A(N4588));
NAND2X1 NAND2_1387 (.Y(N4629),.A(N4569),.B(N4506));
INVX1 NOT1_1388 (.Y(N4630),.A(N4569));
INVX1 NOT1_1389 (.Y(N4635),.A(N4576));
NAND2X1 NAND2_1390 (.Y(N4636),.A(N4576),.B(N4291));
INVX1 NOT1_1391 (.Y(N4640),.A(N4581));
NAND2X1 NAND2_1392 (.Y(N4641),.A(N4581),.B(N4461));
INVX1 NOT1_1393 (.Y(N4642),.A(N4584));
NAND2X1 NAND2_1394 (.Y(N4643),.A(N4584),.B(N4462));
NOR2X1 NOR2_1395 (.Y(N4644),.A(N4608),.B(N4563));
AND2X1 AND2_1396 (.Y(N4647),.A(N4559),.B(N2128));
AND2X1 AND2_1397 (.Y(N4650),.A(N4559),.B(N2743));
BUFX1 BUFF1_1398 (.Y(N4656),.A(N4549));
BUFX1 BUFF1_1399 (.Y(N4659),.A(N4549));
BUFX1 BUFF1_1400 (.Y(N4664),.A(N4564));
AND2X1 AND2_1401 (.Y(N4667),.A(N4587),.B(N4628));
NAND2X1 NAND2_1402 (.Y(N4668),.A(N4413),.B(N4630));
INVX1 NOT1_1403 (.Y(N4669),.A(N4616));
NAND2X1 NAND2_1404 (.Y(N4670),.A(N4616),.B(N4239));
INVX1 NOT1_1405 (.Y(N4673),.A(N4619));
NAND2X1 NAND2_1406 (.Y(N4674),.A(N4619),.B(N4507));
NAND2X1 NAND2_1407 (.Y(N4675),.A(N4186),.B(N4635));
INVX1 NOT1_1408 (.Y(N4676),.A(N4623));
NAND2X1 NAND2_1409 (.Y(N4677),.A(N4623),.B(N4558));
NAND2X1 NAND2_1410 (.Y(N4678),.A(N4365),.B(N4640));
NAND2X1 NAND2_1411 (.Y(N4679),.A(N4368),.B(N4642));
INVX1 NOT1_1412 (.Y(N4687),.A(N4613));
NAND2X1 NAND2_1413 (.Y(N4688),.A(N4613),.B(N4568));
BUFX1 BUFF1_1414 (.Y(N4691),.A(N4593));
BUFX1 BUFF1_1415 (.Y(N4694),.A(N4593));
BUFX1 BUFF1_1416 (.Y(N4697),.A(N4599));
BUFX1 BUFF1_1417 (.Y(N4700),.A(N4599));
NAND2X1 NAND2_1418 (.Y(N4704),.A(N4629),.B(N4668));
NAND2X1 NAND2_1419 (.Y(N4705),.A(N4139),.B(N4669));
INVX1 NOT1_1420 (.Y(N4706),.A(N4656));
INVX1 NOT1_1421 (.Y(N4707),.A(N4659));
NAND2X1 NAND2_1422 (.Y(N4708),.A(N4435),.B(N4673));
NAND2X1 NAND2_1423 (.Y(N4711),.A(N4675),.B(N4636));
NAND2X1 NAND2_1424 (.Y(N4716),.A(N4493),.B(N4676));
NAND2X1 NAND2_1425 (.Y(N4717),.A(N4678),.B(N4641));
NAND2X1 NAND2_1426 (.Y(N4721),.A(N4679),.B(N4643));
BUFX1 BUFF1_1427 (.Y(N4722),.A(N4644));
INVX1 NOT1_1428 (.Y(N4726),.A(N4664));
OR2X1 OR_tmp466 (.Y(ttmp466),.A(N4650),.B(N4350));
OR2X1 OR_tmp467 (.Y(N4727),.A(N4647),.B(ttmp466));
OR2X1 OR_tmp468 (.Y(ttmp468),.A(N4650),.B(N4350));
NOR2X1 NOR_tmp469 (.Y(N4730),.A(N4647),.B(ttmp468));
NAND2X1 NAND2_1431 (.Y(N4733),.A(N4479),.B(N4687));
NAND2X1 NAND2_1432 (.Y(N4740),.A(N4705),.B(N4670));
NAND2X1 NAND2_1433 (.Y(N4743),.A(N4708),.B(N4674));
INVX1 NOT1_1434 (.Y(N4747),.A(N4691));
NAND2X1 NAND2_1435 (.Y(N4748),.A(N4691),.B(N4596));
INVX1 NOT1_1436 (.Y(N4749),.A(N4694));
NAND2X1 NAND2_1437 (.Y(N4750),.A(N4694),.B(N4597));
INVX1 NOT1_1438 (.Y(N4753),.A(N4697));
NAND2X1 NAND2_1439 (.Y(N4754),.A(N4697),.B(N4602));
INVX1 NOT1_1440 (.Y(N4755),.A(N4700));
NAND2X1 NAND2_1441 (.Y(N4756),.A(N4700),.B(N4603));
NAND2X1 NAND2_1442 (.Y(N4757),.A(N4716),.B(N4677));
NAND2X1 NAND2_1443 (.Y(N4769),.A(N4733),.B(N4688));
AND2X1 AND2_1444 (.Y(N4772),.A(N330),.B(N4704));
INVX1 NOT1_1445 (.Y(N4775),.A(N4721));
INVX1 NOT1_1446 (.Y(N4778),.A(N4730));
NAND2X1 NAND2_1447 (.Y(N4786),.A(N4531),.B(N4747));
NAND2X1 NAND2_1448 (.Y(N4787),.A(N4534),.B(N4749));
NAND2X1 NAND2_1449 (.Y(N4788),.A(N4537),.B(N4753));
NAND2X1 NAND2_1450 (.Y(N4789),.A(N4540),.B(N4755));
AND2X1 AND2_1451 (.Y(N4794),.A(N4711),.B(N2124));
AND2X1 AND2_1452 (.Y(N4797),.A(N4711),.B(N2735));
AND2X1 AND2_1453 (.Y(N4800),.A(N4717),.B(N2127));
BUFX1 BUFF1_1454 (.Y(N4805),.A(N4722));
AND2X1 AND2_1455 (.Y(N4808),.A(N4717),.B(N4468));
BUFX1 BUFF1_1456 (.Y(N4812),.A(N4727));
AND2X1 AND2_1457 (.Y(N4815),.A(N4727),.B(N4778));
INVX1 NOT1_1458 (.Y(N4816),.A(N4769));
INVX1 NOT1_1459 (.Y(N4817),.A(N4772));
NAND2X1 NAND2_1460 (.Y(N4818),.A(N4786),.B(N4748));
NAND2X1 NAND2_1461 (.Y(N4822),.A(N4787),.B(N4750));
NAND2X1 NAND2_1462 (.Y(N4823),.A(N4788),.B(N4754));
NAND2X1 NAND2_1463 (.Y(N4826),.A(N4789),.B(N4756));
NAND2X1 NAND2_1464 (.Y(N4829),.A(N4775),.B(N4726));
INVX1 NOT1_1465 (.Y(N4830),.A(N4775));
AND2X1 AND2_1466 (.Y(N4831),.A(N4743),.B(N2122));
AND2X1 AND2_1467 (.Y(N4838),.A(N4757),.B(N2126));
BUFX1 BUFF1_1468 (.Y(N4844),.A(N4740));
BUFX1 BUFF1_1469 (.Y(N4847),.A(N4740));
BUFX1 BUFF1_1470 (.Y(N4850),.A(N4743));
BUFX1 BUFF1_1471 (.Y(N4854),.A(N4757));
NAND2X1 NAND2_1472 (.Y(N4859),.A(N4772),.B(N4816));
NAND2X1 NAND2_1473 (.Y(N4860),.A(N4769),.B(N4817));
INVX1 NOT1_1474 (.Y(N4868),.A(N4826));
INVX1 NOT1_1475 (.Y(N4870),.A(N4805));
INVX1 NOT1_1476 (.Y(N4872),.A(N4808));
NAND2X1 NAND2_1477 (.Y(N4873),.A(N4664),.B(N4830));
OR2X1 OR_tmp470 (.Y(ttmp470),.A(N4797),.B(N4341));
OR2X1 OR_tmp471 (.Y(N4876),.A(N4794),.B(ttmp470));
OR2X1 OR_tmp472 (.Y(ttmp472),.A(N4797),.B(N4341));
NOR2X1 NOR_tmp473 (.Y(N4880),.A(N4794),.B(ttmp472));
INVX1 NOT1_1480 (.Y(N4885),.A(N4812));
INVX1 NOT1_1481 (.Y(N4889),.A(N4822));
NAND2X1 NAND2_1482 (.Y(N4895),.A(N4859),.B(N4860));
INVX1 NOT1_1483 (.Y(N4896),.A(N4844));
NAND2X1 NAND2_1484 (.Y(N4897),.A(N4844),.B(N4706));
INVX1 NOT1_1485 (.Y(N4898),.A(N4847));
NAND2X1 NAND2_1486 (.Y(N4899),.A(N4847),.B(N4707));
NOR2X1 NOR2_1487 (.Y(N4900),.A(N4868),.B(N4564));
AND2X1 AND_tmp474 (.Y(ttmp474),.A(N4823),.B(N4564));
AND2X1 AND_tmp475 (.Y(ttmp475),.A(N4717),.B(ttmp474));
AND2X1 AND_tmp476 (.Y(N4901),.A(N4757),.B(ttmp475));
INVX1 NOT1_1489 (.Y(N4902),.A(N4850));
INVX1 NOT1_1490 (.Y(N4904),.A(N4854));
NAND2X1 NAND2_1491 (.Y(N4905),.A(N4854),.B(N4872));
NAND2X1 NAND2_1492 (.Y(N4906),.A(N4873),.B(N4829));
AND2X1 AND2_1493 (.Y(N4907),.A(N4818),.B(N2123));
AND2X1 AND2_1494 (.Y(N4913),.A(N4823),.B(N2125));
AND2X1 AND2_1495 (.Y(N4916),.A(N4818),.B(N4644));
INVX1 NOT1_1496 (.Y(N4920),.A(N4880));
AND2X1 AND2_1497 (.Y(N4921),.A(N4895),.B(N2184));
NAND2X1 NAND2_1498 (.Y(N4924),.A(N4656),.B(N4896));
NAND2X1 NAND2_1499 (.Y(N4925),.A(N4659),.B(N4898));
OR2X1 OR2_1500 (.Y(N4926),.A(N4900),.B(N4901));
NAND2X1 NAND2_1501 (.Y(N4928),.A(N4889),.B(N4870));
INVX1 NOT1_1502 (.Y(N4929),.A(N4889));
NAND2X1 NAND2_1503 (.Y(N4930),.A(N4808),.B(N4904));
INVX1 NOT1_1504 (.Y(N4931),.A(N4906));
BUFX1 BUFF1_1505 (.Y(N4937),.A(N4876));
BUFX1 BUFF1_1506 (.Y(N4940),.A(N4876));
AND2X1 AND2_1507 (.Y(N4944),.A(N4876),.B(N4920));
NAND2X1 NAND2_1508 (.Y(N4946),.A(N4924),.B(N4897));
NAND2X1 NAND2_1509 (.Y(N4949),.A(N4925),.B(N4899));
NAND2X1 NAND2_1510 (.Y(N4950),.A(N4916),.B(N4902));
INVX1 NOT1_1511 (.Y(N4951),.A(N4916));
NAND2X1 NAND2_1512 (.Y(N4952),.A(N4805),.B(N4929));
NAND2X1 NAND2_1513 (.Y(N4953),.A(N4930),.B(N4905));
AND2X1 AND2_1514 (.Y(N4954),.A(N4926),.B(N2737));
AND2X1 AND2_1515 (.Y(N4957),.A(N4931),.B(N2741));
OR2X1 OR_tmp477 (.Y(ttmp477),.A(N2483),.B(N4921));
OR2X1 OR_tmp478 (.Y(N4964),.A(N2764),.B(ttmp477));
OR2X1 OR_tmp479 (.Y(ttmp479),.A(N2483),.B(N4921));
NOR2X1 NOR_tmp480 (.Y(N4965),.A(N2764),.B(ttmp479));
INVX1 NOT1_1518 (.Y(N4968),.A(N4949));
NAND2X1 NAND2_1519 (.Y(N4969),.A(N4850),.B(N4951));
NAND2X1 NAND2_1520 (.Y(N4970),.A(N4952),.B(N4928));
AND2X1 AND2_1521 (.Y(N4973),.A(N4953),.B(N2739));
INVX1 NOT1_1522 (.Y(N4978),.A(N4937));
INVX1 NOT1_1523 (.Y(N4979),.A(N4940));
INVX1 NOT1_1524 (.Y(N4980),.A(N4965));
NOR2X1 NOR2_1525 (.Y(N4981),.A(N4968),.B(N4722));
AND2X1 AND_tmp481 (.Y(ttmp481),.A(N4946),.B(N4722));
AND2X1 AND_tmp482 (.Y(ttmp482),.A(N4818),.B(ttmp481));
AND2X1 AND_tmp483 (.Y(N4982),.A(N4743),.B(ttmp482));
NAND2X1 NAND2_1527 (.Y(N4983),.A(N4950),.B(N4969));
INVX1 NOT1_1528 (.Y(N4984),.A(N4970));
AND2X1 AND2_1529 (.Y(N4985),.A(N4946),.B(N2121));
OR2X1 OR_tmp484 (.Y(ttmp484),.A(N4954),.B(N4344));
OR2X1 OR_tmp485 (.Y(N4988),.A(N4913),.B(ttmp484));
OR2X1 OR_tmp486 (.Y(ttmp486),.A(N4954),.B(N4344));
NOR2X1 NOR_tmp487 (.Y(N4991),.A(N4913),.B(ttmp486));
OR2X1 OR_tmp488 (.Y(ttmp488),.A(N4957),.B(N4347));
OR2X1 OR_tmp489 (.Y(N4996),.A(N4800),.B(ttmp488));
OR2X1 OR_tmp490 (.Y(ttmp490),.A(N4957),.B(N4347));
NOR2X1 NOR_tmp491 (.Y(N4999),.A(N4800),.B(ttmp490));
AND2X1 AND2_1534 (.Y(N5002),.A(N4964),.B(N4980));
OR2X1 OR2_1535 (.Y(N5007),.A(N4981),.B(N4982));
AND2X1 AND2_1536 (.Y(N5010),.A(N4983),.B(N2731));
AND2X1 AND2_1537 (.Y(N5013),.A(N4984),.B(N2733));
OR2X1 OR_tmp492 (.Y(ttmp492),.A(N4973),.B(N4475));
OR2X1 OR_tmp493 (.Y(N5018),.A(N4838),.B(ttmp492));
OR2X1 OR_tmp494 (.Y(ttmp494),.A(N4973),.B(N4475));
NOR2X1 NOR_tmp495 (.Y(N5021),.A(N4838),.B(ttmp494));
INVX1 NOT1_1540 (.Y(N5026),.A(N4991));
INVX1 NOT1_1541 (.Y(N5029),.A(N4999));
AND2X1 AND2_1542 (.Y(N5030),.A(N5007),.B(N2729));
BUFX1 BUFF1_1543 (.Y(N5039),.A(N4996));
BUFX1 BUFF1_1544 (.Y(N5042),.A(N4988));
AND2X1 AND2_1545 (.Y(N5045),.A(N4988),.B(N5026));
INVX1 NOT1_1546 (.Y(N5046),.A(N5021));
AND2X1 AND2_1547 (.Y(N5047),.A(N4996),.B(N5029));
OR2X1 OR_tmp496 (.Y(ttmp496),.A(N5010),.B(N4472));
OR2X1 OR_tmp497 (.Y(N5050),.A(N4831),.B(ttmp496));
OR2X1 OR_tmp498 (.Y(ttmp498),.A(N5010),.B(N4472));
NOR2X1 NOR_tmp499 (.Y(N5055),.A(N4831),.B(ttmp498));
OR2X1 OR_tmp500 (.Y(ttmp500),.A(N5013),.B(N4338));
OR2X1 OR_tmp501 (.Y(N5058),.A(N4907),.B(ttmp500));
OR2X1 OR_tmp502 (.Y(ttmp502),.A(N5013),.B(N4338));
NOR2X1 NOR_tmp503 (.Y(N5061),.A(N4907),.B(ttmp502));
AND2X1 AND_tmp504 (.Y(ttmp504),.A(N5021),.B(N4991));
AND2X1 AND_tmp505 (.Y(ttmp505),.A(N4730),.B(ttmp504));
AND2X1 AND_tmp506 (.Y(N5066),.A(N4999),.B(ttmp505));
BUFX1 BUFF1_1553 (.Y(N5070),.A(N5018));
AND2X1 AND2_1554 (.Y(N5078),.A(N5018),.B(N5046));
OR2X1 OR_tmp507 (.Y(ttmp507),.A(N5030),.B(N4335));
OR2X1 OR_tmp508 (.Y(N5080),.A(N4985),.B(ttmp507));
OR2X1 OR_tmp509 (.Y(ttmp509),.A(N5030),.B(N4335));
NOR2X1 NOR_tmp510 (.Y(N5085),.A(N4985),.B(ttmp509));
NAND2X1 NAND2_1557 (.Y(N5094),.A(N5039),.B(N4885));
INVX1 NOT1_1558 (.Y(N5095),.A(N5039));
INVX1 NOT1_1559 (.Y(N5097),.A(N5042));
AND2X1 AND2_1560 (.Y(N5102),.A(N5050),.B(N5050));
INVX1 NOT1_1561 (.Y(N5103),.A(N5061));
NAND2X1 NAND2_1562 (.Y(N5108),.A(N4812),.B(N5095));
INVX1 NOT1_1563 (.Y(N5109),.A(N5070));
NAND2X1 NAND2_1564 (.Y(N5110),.A(N5070),.B(N5097));
BUFX1 BUFF1_1565 (.Y(N5111),.A(N5058));
AND2X1 AND2_1566 (.Y(N5114),.A(N5050),.B(N1461));
BUFX1 BUFF1_1567 (.Y(N5117),.A(N5050));
AND2X1 AND2_1568 (.Y(N5120),.A(N5080),.B(N5080));
AND2X1 AND2_1569 (.Y(N5121),.A(N5058),.B(N5103));
NAND2X1 NAND2_1570 (.Y(N5122),.A(N5094),.B(N5108));
NAND2X1 NAND2_1571 (.Y(N5125),.A(N5042),.B(N5109));
AND2X1 AND2_1572 (.Y(N5128),.A(N1461),.B(N5080));
AND2X1 AND_tmp511 (.Y(ttmp511),.A(N5055),.B(N5085));
AND2X1 AND_tmp512 (.Y(ttmp512),.A(N4880),.B(ttmp511));
AND2X1 AND_tmp513 (.Y(N5133),.A(N5061),.B(ttmp512));
AND2X1 AND_tmp514 (.Y(ttmp514),.A(N5085),.B(N1464));
AND2X1 AND_tmp515 (.Y(N5136),.A(N5055),.B(ttmp514));
BUFX1 BUFF1_1575 (.Y(N5139),.A(N5080));
NAND2X1 NAND2_1576 (.Y(N5145),.A(N5125),.B(N5110));
BUFX1 BUFF1_1577 (.Y(N5151),.A(N5111));
BUFX1 BUFF1_1578 (.Y(N5154),.A(N5111));
INVX1 NOT1_1579 (.Y(N5159),.A(N5117));
BUFX1 BUFF1_1580 (.Y(N5160),.A(N5114));
BUFX1 BUFF1_1581 (.Y(N5163),.A(N5114));
AND2X1 AND2_1582 (.Y(N5166),.A(N5066),.B(N5133));
AND2X1 AND2_1583 (.Y(N5173),.A(N5066),.B(N5133));
BUFX1 BUFF1_1584 (.Y(N5174),.A(N5122));
BUFX1 BUFF1_1585 (.Y(N5177),.A(N5122));
INVX1 NOT1_1586 (.Y(N5182),.A(N5139));
NAND2X1 NAND2_1587 (.Y(N5183),.A(N5139),.B(N5159));
BUFX1 BUFF1_1588 (.Y(N5184),.A(N5128));
BUFX1 BUFF1_1589 (.Y(N5188),.A(N5128));
INVX1 NOT1_1590 (.Y(N5192),.A(N5166));
NOR2X1 NOR2_1591 (.Y(N5193),.A(N5136),.B(N5173));
NAND2X1 NAND2_1592 (.Y(N5196),.A(N5151),.B(N4978));
INVX1 NOT1_1593 (.Y(N5197),.A(N5151));
NAND2X1 NAND2_1594 (.Y(N5198),.A(N5154),.B(N4979));
INVX1 NOT1_1595 (.Y(N5199),.A(N5154));
INVX1 NOT1_1596 (.Y(N5201),.A(N5160));
INVX1 NOT1_1597 (.Y(N5203),.A(N5163));
BUFX1 BUFF1_1598 (.Y(N5205),.A(N5145));
BUFX1 BUFF1_1599 (.Y(N5209),.A(N5145));
NAND2X1 NAND2_1600 (.Y(N5212),.A(N5117),.B(N5182));
AND2X1 AND2_1601 (.Y(N5215),.A(N213),.B(N5193));
INVX1 NOT1_1602 (.Y(N5217),.A(N5174));
INVX1 NOT1_1603 (.Y(N5219),.A(N5177));
NAND2X1 NAND2_1604 (.Y(N5220),.A(N4937),.B(N5197));
NAND2X1 NAND2_1605 (.Y(N5221),.A(N4940),.B(N5199));
INVX1 NOT1_1606 (.Y(N5222),.A(N5184));
NAND2X1 NAND2_1607 (.Y(N5223),.A(N5184),.B(N5201));
NAND2X1 NAND2_1608 (.Y(N5224),.A(N5188),.B(N5203));
INVX1 NOT1_1609 (.Y(N5225),.A(N5188));
NAND2X1 NAND2_1610 (.Y(N5228),.A(N5183),.B(N5212));
INVX1 NOT1_1611 (.Y(N5231),.A(N5215));
NAND2X1 NAND2_1612 (.Y(N5232),.A(N5205),.B(N5217));
INVX1 NOT1_1613 (.Y(N5233),.A(N5205));
NAND2X1 NAND2_1614 (.Y(N5234),.A(N5209),.B(N5219));
INVX1 NOT1_1615 (.Y(N5235),.A(N5209));
NAND2X1 NAND2_1616 (.Y(N5236),.A(N5196),.B(N5220));
NAND2X1 NAND2_1617 (.Y(N5240),.A(N5198),.B(N5221));
NAND2X1 NAND2_1618 (.Y(N5242),.A(N5160),.B(N5222));
NAND2X1 NAND2_1619 (.Y(N5243),.A(N5163),.B(N5225));
NAND2X1 NAND2_1620 (.Y(N5245),.A(N5174),.B(N5233));
NAND2X1 NAND2_1621 (.Y(N5246),.A(N5177),.B(N5235));
INVX1 NOT1_1622 (.Y(N5250),.A(N5240));
INVX1 NOT1_1623 (.Y(N5253),.A(N5228));
NAND2X1 NAND2_1624 (.Y(N5254),.A(N5242),.B(N5223));
NAND2X1 NAND2_1625 (.Y(N5257),.A(N5243),.B(N5224));
NAND2X1 NAND2_1626 (.Y(N5258),.A(N5232),.B(N5245));
NAND2X1 NAND2_1627 (.Y(N5261),.A(N5234),.B(N5246));
INVX1 NOT1_1628 (.Y(N5266),.A(N5257));
BUFX1 BUFF1_1629 (.Y(N5269),.A(N5236));
AND2X1 AND_tmp516 (.Y(ttmp516),.A(N5254),.B(N2307));
AND2X1 AND_tmp517 (.Y(N5277),.A(N5236),.B(ttmp516));
AND2X1 AND_tmp518 (.Y(ttmp518),.A(N5254),.B(N2310));
AND2X1 AND_tmp519 (.Y(N5278),.A(N5250),.B(ttmp518));
INVX1 NOT1_1632 (.Y(N5279),.A(N5261));
INVX1 NOT1_1633 (.Y(N5283),.A(N5269));
NAND2X1 NAND2_1634 (.Y(N5284),.A(N5269),.B(N5253));
AND2X1 AND_tmp520 (.Y(ttmp520),.A(N5266),.B(N2310));
AND2X1 AND_tmp521 (.Y(N5285),.A(N5236),.B(ttmp520));
AND2X1 AND_tmp522 (.Y(ttmp522),.A(N5266),.B(N2307));
AND2X1 AND_tmp523 (.Y(N5286),.A(N5250),.B(ttmp522));
BUFX1 BUFF1_1637 (.Y(N5289),.A(N5258));
BUFX1 BUFF1_1638 (.Y(N5292),.A(N5258));
NAND2X1 NAND2_1639 (.Y(N5295),.A(N5228),.B(N5283));
OR2X1 OR_tmp524 (.Y(ttmp524),.A(N5278),.B(N5286));
OR2X1 OR_tmp525 (.Y(ttmp525),.A(N5277),.B(ttmp524));
OR2X1 OR_tmp526 (.Y(N5298),.A(N5285),.B(ttmp525));
BUFX1 BUFF1_1641 (.Y(N5303),.A(N5279));
BUFX1 BUFF1_1642 (.Y(N5306),.A(N5279));
NAND2X1 NAND2_1643 (.Y(N5309),.A(N5295),.B(N5284));
INVX1 NOT1_1644 (.Y(N5312),.A(N5292));
INVX1 NOT1_1645 (.Y(N5313),.A(N5289));
INVX1 NOT1_1646 (.Y(N5322),.A(N5306));
INVX1 NOT1_1647 (.Y(N5323),.A(N5303));
BUFX1 BUFF1_1648 (.Y(N5324),.A(N5298));
BUFX1 BUFF1_1649 (.Y(N5327),.A(N5298));
BUFX1 BUFF1_1650 (.Y(N5332),.A(N5309));
BUFX1 BUFF1_1651 (.Y(N5335),.A(N5309));
NAND2X1 NAND2_1652 (.Y(N5340),.A(N5324),.B(N5323));
NAND2X1 NAND2_1653 (.Y(N5341),.A(N5327),.B(N5322));
INVX1 NOT1_1654 (.Y(N5344),.A(N5327));
INVX1 NOT1_1655 (.Y(N5345),.A(N5324));
NAND2X1 NAND2_1656 (.Y(N5348),.A(N5332),.B(N5313));
NAND2X1 NAND2_1657 (.Y(N5349),.A(N5335),.B(N5312));
NAND2X1 NAND2_1658 (.Y(N5350),.A(N5303),.B(N5345));
NAND2X1 NAND2_1659 (.Y(N5351),.A(N5306),.B(N5344));
INVX1 NOT1_1660 (.Y(N5352),.A(N5335));
INVX1 NOT1_1661 (.Y(N5353),.A(N5332));
NAND2X1 NAND2_1662 (.Y(N5354),.A(N5289),.B(N5353));
NAND2X1 NAND2_1663 (.Y(N5355),.A(N5292),.B(N5352));
NAND2X1 NAND2_1664 (.Y(N5356),.A(N5350),.B(N5340));
NAND2X1 NAND2_1665 (.Y(N5357),.A(N5351),.B(N5341));
NAND2X1 NAND2_1666 (.Y(N5358),.A(N5348),.B(N5354));
NAND2X1 NAND2_1667 (.Y(N5359),.A(N5349),.B(N5355));
AND2X1 AND2_1668 (.Y(N5360),.A(N5356),.B(N5357));
NAND2X1 NAND2_1669 (.Y(N5361),.A(N5358),.B(N5359));
endmodule 